PK   c��T�t��`  �    cirkitFile.json���q&�*ݿXDF^��?�a���B�p7 l��"�"��b�#��e�&s��ɽ*�VeV|AK<�u�2���TdFTfğ^���m~�0�{??������wo_�@�����?���V�|����=�����߿��O鿛�������~��9��϶�F�vj,�i�l5̴R��zP/~��/�S 6�@l\
�A�1p)������,��zpl\
���1p)�������Z6.�б1p)D�w�l�U�}%�%�DD�w�l�a�ID|��&Q�&�DD����?���������j���Sm��jm��fi��?�n�B�`�&|�K|��&Qt7r����������r?�{ӿ��?���r�������$"
�g��( ^��|�&QX��pL��|�����M"���6����mf��(�>�M"��o��$b\���l��ID|��&Q R|�k�{g6����;�$"
�０8��)�*��v�oM@n߅�g��(�.�MB=X�g��(�.�M"��p6������$"
@����-߅�I��:`��o-+����>��A�‸�}���l6	��sEv
�";��w|��&Q��?�DDa8oI����r��~�ϟ�}�r�p	�r�_�b��(�i6�����g��(����z��=<�DD���l߇g$����_;�\�c��X��>���inô��y�/`H�J�@bXH(�C	1�Ck��ȭ{N̅��yi�ֹ�z56���F�=�!x���(��䦱j�85КOnPF3l\��}Q/7���d!�3�a�C��b���a��!Vv+;(:¢�[7��<VvPt���ڃ��#�����76:����~CC���ȵ�C��m+��{���m�r�Z��[�ܡ��N=tX�uX�A�]:�:�p�����#0�tT,?h0C`|Ɨ����B������x�������`��,>�KW��9X|Ɨ.S��t���/]��`�_���8���#0���/�e�{��/��m��L���_���/�R��`�_�_�8|��#0�t3,?p���G`|�NX~������ҍ:�����񥻀`���,>�K����/X|Ɨ�_��_���/������6�m}A�~�'���/��Xgl��06-9�'e�n$�Y<]8t���`�YKw���G=X|Ɨn7���z���/���}"}$�p�c�Q���`���,>�K����G=X|�w[ "�,��$�M�nW�AS�S\�ɀ�&,>�K���MX|Ɨ�L`�g�����`���,>�K�=���/X|��o+��zj���w���]��5����i0�R�+n�Xp��;-*�s,k��X��<�<�ɂ�&����/���4a�_����S��zC`��������'�A�CcC�ͳo:\�6h��6L3�L0Yp���G`|�� I��<8U��'.,{��S\�xˁ�-,>��w��ʄ�"\`уC5,>�K�����[X|Ɨ�czJ�}�1W��D��

�
�
��ˁc.�����/U��sa�_���8���#0�TQ,?p���G`|�"V~��	����RG��������`���,>:�Wݪ��۾4�`<}]|�r��jh��u���fU����ĕ��U�k�V���VN_�5�u����L�#��]zen�.:�Xo�j�֖����}�5,���9=ڲ�|_��������dMk�3_��1a�|��g�j�3�u�D�v>����u�+-���fq����6���m���0�y����w��;��b=zo�)*_�Zm��jS�h�z4�m�z��n��o{�W�v>s�������X����E���Y���xby�Uӭ����:f�x�c=��>���U��J�ŊL.ݤN?��Ld-�j�3��.О�^�}S�x����M��]�z<��8���Z"��g.�Y�����:k�S;���y�b�y<fh虡�gڟg�_`�_`�_`�_`�_`�_`�_�&������7L���8��}@����<���g��-��i�/O�|yZ���2_������L��1�w�t���:��uL���u(-������ɅJ?OW�˿N�﮹�mtA����O��/>�q�	!��𝎆���UEO�jrS������49��-p(�9�~�kd�)�ץz����&�0.9�+�\Y���[�z��?�&�0.�)��!��������C59����U�Ȭ&���:īx���jr�q����YM��u�]/�������k_�|��w�w��``�Բ���Q�S�8zK��Y�:�U�y�tZ���g�t�WW�jr��= =�Ň��쉌?eWް����,������" q���A�Q�g��3n==��9����� Z�ݰ,��=�E~����n==��3,�G]�Oh���*o�[O�E~���Q��Z����	�Ӄh���²x�1���Y����� Z�'��,�m>�E~�r==��,�t����"7RӀ��D����ţ�'����������"�ŚV��� G4����n��� �4��,�G�Oh���)�]O�E~���Q[�Z��B�B���B���n��'�����~B����ţ�'���ݔw1�����%�2_bj����Ӡ�i����� ��b�i ������@<?�U�羞Ġ��;����0��T^F����0·齲3�����Ұ�Qy!���48��y��(�� 8/���),�A��z���ഞ�X.e�C���N	f��N\��8%�f��,�E�W<!upJЀS�l	�"�YT�:�L��S��d�H`	̢���dJ}�}�p�Ĳ��UG�R�8%�*�Z_ꏩ1p
+u-���8�g�9��ڶ��&�#ÊG]��25N�p�m��pi�S���)7�xԵ2Sc�����v+=��&gj�rÊG�ըOh�r3������25x���)�pp �O�p�̀Sn���
S��\..��x�ի�7 ��Yp��"�Y$0�*�pB���g��,�E����'���Yp��"�Y$0�*�qB���g��,�E���>&'���=�.>�>�.?��Y~΂�p��c�H`	̢�6�aJ�I��L�E�H`յ�S��l�g��,�E���-��Rg�,8��f��,�Eu�Ŕ:8�d�i$6�f��,�k�2��8w���6�f��,�k�7�����ݰY$0�fQ�m�NH��q���E�H`U��������ݰY$0�fQ][J2���8p��"�Y$0��ڙ�)ut�xt�x@�xtyp���s7��q�܍c��r�SPX�X<��c��1p�ǁ�>l	�"�YTy��R�}8��Z�{�-܍�ţ�f�'4�9pΈ�"�Y$0�*oy]/u�yp��+�{�-ހ�ţ��'4�7yp���"�Y$0�*oB��|��.,���w����|��i��J�f��X����yj�O�&�{�u�����z�h�~����T�����E���^M��z]4}��u�����E��[^����v��s��ϴ���}��}���`F5G�A>��m��u���Sl��~ו���Oa���$5�хS�ye�@�i�=��Ӌ��?�׋j'�7\���im�yR-�n�ź;O/����I7�07a	q5��jz�l�n����@흧M��RZ�~�ӽ���cד�Y��v��iR��}������s�U�Y�E���n�z����l�M��]l�G]3��6֌�B77�Ҽ�y��|�����O�ޘ0X��t4�o�t�wd���{z/����h�q3�fj繱��7�8����^5�yz�t������H5Ɨ-�S���7��	C�[z���6
{�_*�K���a@!�F�8Σ�B4L!�?s�I:�A׎�{�9�5�q]\=���i0�R|}�i4]	��P��+����ߢ�c��9�Y�(�<��q����ĵȺ��!FD䜏��܍��JА�<�k:�ZN(�	e]�kJ;�w/C���(�;��f�l4A���{M�����h��;T4}S_4}O_4}K_4}?�,��NM�'��ef�5;���	'��3-�N8Y6��M!�Ω!���i��ѸK�ŹiGko{Y2�NP��Y�`�q��qz�1���<���&?wzw{Gԛ!�No�(F�}t�Au��ȵÃ��vEO��=yo7X�佌fѓ�V��'�m4�����=yo�Q��v��E�y߁�Ѭ���Ѭ���SuѣY�Y�g߅a�х����*X������;���体���佳V������$e�u_�[/s.�P<��0��Ѕ8y���u��}܂x?ء��l!���o!����ߺ���%�L������@�Ԏ]g��/�t|��}���?�oB�&h���A9�ۻ��E��^b�h:����+�����<x׶��K�nf�tdMcf2�6��t/�_4}��Eޛn;=�8��M||�v��0-�`ؙ��@n6B���"$�d�ʄ��T�L�|��������ͻ�/~����%R�Ë��.���9�P�:�K2�D�� ��Y1�@�.�W"!���D B*��0�@�T�qc���� Ri��A"�.�e���ym�ۆ�m�9n%uɱ�0�|7��7����A�`��`EI���Ҳ�̇̉�(][�'J��1�����q�k;m&�����q��(J�ƽ_�a~\��8�ҵ}(̏k�VE��`�	��5l;��t�
�a~���8�ҵ�.��K�������Q���@�`~�����������P�L����Q���@�`~���8�ҵ>̏[�GQ�V)a���qIq��0?��t���ۏۋ����	��m�����Q��uD1k���q��(J�� L0?���̏����կ r�}��}ބ�q��(J�j] L0?�`�q�k5$&����8�ҵ�̏{�ߣ�>?��?�g�6Wy��7��,�zX���hk]�#W	����/�uq8U�\%��&V�֥�1~`]`#�+�*P��b�p�@�J`%�q$"�ub�$��V��.��
����h?�.�����.F9V�>K�zX��S�U+�`U�r�p�@�J`%��L�L`�� ��hIm:�,#[�H�dВ�tF[F��ɠ%�鬹�le�/�$�6�����L&��dЦ��2����DВ�t�AF�2��Z�A��b��V&AK2hӝ��Dd"hIm�##ۭH�UA&,�D����˴L\&��dЦ�J2����DВ�t�JF�2q�Z�A����V&.AK2h�8���e"hIm��'#[��L-ɠMwed+���%��n��le�2�$�6����L\&��dЪ���H��|-A�W�}7_׽Gw���6�">���Mw�ed+���%����le�2�$�6�����iE��2q���ˌL\&��dЦ��2����DВ�Tc@F�2q�Z�A�j%��v+��wAK�hB��ˌL\&��dЦ�2����DВ�T�CD�V&.AK2hS-���e"hI��i����L\&�6�C	�լ;m�d+�m�E�jDЦ52��I&t�L&.�2q����DВ�T3HF�2q�Z�A�j��V�{�Z�A��.�d����B�2�����eV&.AK2hSM-�:��"hi-@2q����D��6Z~��d�2'���%��V��le�2�$�6՜Xyo�"e+���M��d�V�ʇP������eN&.AK2hS-C���e"hIm��(#[��L-ɠM�%ed+���%��F��l���2�$�6�����L\&��dЦ��2����D�R�g�Qm׵����R�m��,M;y��MS�}��N&�Tvj�VR٩&[Ie��w%���ەTvjeWR٩n]Ie�u%��
ҕTvj>�Z�N��Z2�%��^��.����!�1�n��d.&��R��!0d0F��ٳ��a�x�f-��u��%���^��d0�x��b-���5�]u1V��=���Ŋ�2��r��!s��Q�c�٫=��������uu���a�x�wZ-�/��1�_���]�k�x� y5���d:��6T�W�s�Ɗ��3Ւ�6��Es���.H|2C&`�`|�^G�ڨ����Ԓ�X��X���b�O`���/�+�+++++++�4ƊƊ�Ŋ����Y?�!C2+n1V�b���Xq����-�Xq����w_�a���Xq��⮠;�Au��̭s��jlZ=����z�C�&��;�jVH��[\5��Oq�L���`�0�����z��~Ѯ��{и^� ��&VSj��]h!!M�|^��4���>��Ta��>����v5U��ALou�����*���7���Lx5U��AL�����
���֮^'�'ԫ�5b���f5U��wb�z�Ԟ���
�4���~��T���	��uR{z��*P����v(��
�t�����I�]�j��(k'�T�	��z��kz'YV��ڛ�T���Η�z�H0]���D��$��ZO�l�':�֓E��*ʕI����n��d���%̪;�֓E��3Ự�	}��f��q��"�˜��]����aɳꎽ�d�����D�.�T|B߰Zu�z�H}òh"|vO>�oX"���q=Y��a�4�;:��7,�V�m��,R� �Ot��'��7(�t�_u=Y��ay5�;_��7,�Vݕ��,R� �Ot�'�<�˯Uwʮ'�<�˯��]�!���a������d�����D�.�Z~B߸iB'҄���Τ	J�ɯ�U%8���ZQ������D�.��~B߰�Zu��z�H}[������O����8���ZQ7��v��'|��"�oX~��C}=Y��=괃�$÷ڭ�sB12�5-�_�;U*N(F&�&·�-qtB12�5-�_Ӡ�z$�7m�X�a�5-�_�2�5;�&�7��v�����#�_32�5�$�7��v���P�L~����P|��$÷z,�Q�L~����P|��$÷z��Q�нO������2�5��caK�bd�kF&��W��bd�k"|��
����׌L~��7D�2��D�V�K�#�_32�5˯��M2|��5}��ɯ������D�&��n����ɯ��ڕoHM�ڎ��d����׌L~���מ���SE��m���Խr����2�5+�_C�M2|��j���	���׬L~�7��M2|��'#�_�2�5�$�7��v;9�P�L~����P|��$÷�m�qB1B�Մʫ��	X�ɯYX~���׬L~�7��M2|��&6���׬L~�7��M2|��nC���׬L~�7��M2|�ǶP���׬L~�7��M2|���]���׬L~�7��M2|�ύ���q2�5'�_C�M2|���sG<�bd�kN&���d�&��n����ɯ9���o��d�V�=&O(F&��d�k(�I�o��[=6�(F&��d�k(�I�o��[=vm�(F���P\�62�5˯9����ɯ�>������2D12�5'�_C�M2|��j�a�	���לL~��7���ɯ��v;��P�L~����P|��$÷�m_�/�_�2��+߈�[�o��;��_�2�5/�_C�M2|��Q�����ɯy��ڕo��-�_+��Kkh�u7+�i�Cc�⛞�YL?������^o�J*�������.���5��r�x���a��"*��㋨��/�r�:���a��2�/�z�ڣԒ���^3�Z2�����j�Ί|$3��c�ғ��>�����r�'
����y�~t���+���HC���c)�r��׋j'�7\�HMs���5�Z"��u�X��b�Tps��6vV�鍳�[�qng��X��bQJ��/��Wq��ql���5�3�N};M�`U*�r�%�����ڨ�.�]�-Q���S�M8�RD��]lM]3��6֌�B77�Ҽ�y��\ �"*�X�7&V5�#���k��n�����B�P`/ET�Do�nR���sc��o�q69=,&��j<�RD��p����:�~����Nׄ��-��|�(��XI��Ѩ۱[T0=�k��s�lWG�v���8�5�q]\���i0�R�r)�B,�r)�r���* *��
��<955~��Һ���r�Go9w#]��,Jw�
騈�>�Q;��-C���(�{�huq�M�m���3Q9�ET��������������a|SD�0�)�r�Q9�oʬd��=�o��`��8�)#sh�����fj�,iӧ0)�hqn������?J���<��m�h|�I&�5����ϝ~��s۱�\�S�c����\L&n�Z���g�@*��ݲLz���;��qU�&�bb���H����qt���I�6�aP!�b T��QqGVWD%�K�b/��(��S)���7ϳ�qcl��čYk���3��Џ��ή�ʡ�+�r�&u��;K��F�6�$bh�"Fpcי���6sTD吣Q���7!D�d���A�&�hf}U�
B�"*,��-�r���޵m����Y7YӘ�̠c��� UVD�P.��71 �!��T�ܴ�O���inô��9B���ET4�����2�=|���_���jS?�v��\�RL��9���L�!5��>\�����7{��J��5�� �& �@��I	"�k��DH]6+D B�ـ R�����l� �@��esA"��E���ym�ۆ�m�9n%uͯ`0�|7��7���f~0�`��`E�{:̇̉�(=v��`��q��(J��|1�p�o���5̏�(=v��`��q��(J�1�`~\��8��c'9&��0?���ؑ������q���FL�L
.�����Q���`0�����q��nL0?n`~E鱪>̏[�GQz�N������Q��<c0�r⸤8̏[�GQz�������Q�+cb0�����q��
��O?0?�`~E�R̏;�GQz�x��������	����Q���`0�����q��*!L0?�a~E��̏{�ߣ��2|Ṣ�{4��{ U�J"X�CV�M(W	�$�U=d%!�T�r��J"X�CV�M(W	�$�5�]"r�*�B$ ��D��}��\�J�	H`%�q�""׬"&DXI�z�JO���*��D�����#�*P�XI�z�J)���*��D��3�2��L�%��dЦ��2�����.���d/���DВ�t�\F�2їZ�A�����V&AK2h����Da"hIm�� #[�HL-ɠMw1dd+���%��N��le"2�$�6ݍ���LT&��dЦ;>2d�2�$�6�U���L\&��dЦ;W2��"&�IL&.�2q����DВ�tNF�2q�Z�A�����V&.AK2hӝD���e"hIm�[)#[��L-ɠMwDed+���%�鮫�le�2�$�6�ٕ9�$���%��le�2�$�6ݡ���L\&��dЦ��2�:�(t\Q&.32q����DВ�t7_F�2q�Z�A�j��V&.AK2hS����e"hIm�� #[��L-ɠM�+dd+���%����l�L\&��dЦZ"2����DВ�TEF�2q�Z�A�j���V&.AK2hS��
�$�J&�Y�����e"hIm�$#[��L-ɠM��dd+���%�����le�2�$�6բ���L\&��dЦ�Z"�u2q�Z�A�j���V&.AK2hS�3���e"hIm��&#[��L-ɠM5�dd+���%��v��l��|����˜L\�d�2�$�6�2���L\&��dЦ��2����DВ�T[RF�2q�Z�A�jd�����e"hIm��)#[��L-ɠM5Ked+����2��ZE{�ڮk#A��Z�t�Y�v��������a���S����N5�J*;u�+��Tޮ��S+���Nu�J*;��+��T����S���@Ƌ�^�^��Z2��ZKc�{=Gk�`�x��g���X�^��Z2+��RYKc�{� k�`�x��b-���5�]u1V��=��h+��⽶z�d0V�׼��Ɗ�Z�Ւ�X�^#�Z2+�kwVK�#�X�^�Z2+��UKc�{=�j���u��%����L�d@�Ɗ�Ւ�X�^{�Z2+�k�SKc�{�nj�`��c�؃�+�+�+�+++++++�4ƊƊƊ[��+n1V�b���Xq���c�-([���c�Ɗ;�w+�0V�a��+��BPݼ4s�\c��VO}�㿇���I�������WMu�S\-ӄb��Ga5U�j��a�Nj�hWSj�t}��j�@M�-$$������1]�Ǳ�*P�;�R�NjOaWSj�t}g�j�@M���uR{&��*P� ��{]VSjzgkW�����T��1]�}��*P�;1d�Nj��WSj�t}?�j�@M���:�=�_M�i��J��5�����I�]�j�@M����ZM��dY�Njo6TSj�t}�j���	,IV�a��,2y˓��]�Y���q�2�\�P��-J��������P�LƬ��	}�rf"|v�=�oXڬ�;n=Y��a�3����7,yVݱ��,R߰��߅��O��B��"\O�oXM�����'�K�Uw6�'��7,�&�waG����Ӫ�-דE��QỰ��	}Òj����"�˫��]�����a�����d���e�D�.��}�
,�V�)��,��
,�&�wa�����ת�wדE��_Ựk�	}��	�H:��;�&t(M&��W���bd�kE]�O��_Ự��	}��k՝���"�˯��]�q���a���n��d�����D�&��nA���ɯu�?�oX~M�o��[�V�9�����ɯ��&�I�o�[��bd�kZ&���d�&��n-���ɯi���o��d�V�E�N\�ɯ���o��d�V���N(F&�fd�k(�I�o��[��;�����ɯ��&�I�o�[/�b��}
]������)�_�+lyB12�5#�_C�M2|��j��	���׌L~�7��M2|��R�'#�_32�5�$�7��vk��P�L~����P|��$÷�-�|B12�5#�_C�M2|��j�J�	���׌L~�7��M2|��r����2�5+�_C�M2|��j���	���׬L~�7��M2|��'#�_�2�5�$�7��v;9�P�L~����P|��$÷�m�qB1B�Մʫ��	X�ɯ��F9�����ɯ��&�I�o����bd�kV&���d�&��n����ɯY���o��d�V�m�N(F&�fe�k(�I�o��[���:�����ɯ��&�I�o��h�^1N&��d�k(�I�o��[�v�;�����ɯ��&�I�o�ۺ��bd�kN&���d�&��n����ɯ9���o��d�V��@O(F&��d�k(�I�o��[�vm=��BMp]��������P�L~����P|��$÷��|B12�5'�_C�M2|��j�a�	���לL~�7��M2|����'#�_s2�5�$�7��v[��+���׼L~�7��M2|Gq��k^&��e�k(�I�o��;��_�2�5/�_C�M2|S�_ZC;��Yi�L����4O�b�i���}o�zWR9�]D��v���Y%����ET��Q9l_D�w|����ET;ǗY�x1ֻ����~��9Ԓ9�`�fTstV�#��ئ[א��<���n�m|%�C=Qf��8W�c����t^�&��G�ń�K�C,�^T;龡�"Gj���v��'��vX�;�RD�ˤ��h�������RMo�m�ҍs�8�=�RD��RZ�~�T��k�c���Y��v��iR�R�C,a�ܼh�t�FMw�=��n������l�1�"*�X�b#h�Q��f����1�����l��Q9Ģ�1a����hu]�t�wd���{)�r�%Zx�u�j�v��/}ӎ�i��a1�T�1�"*,�ˀ�H5��9�S|�f�t:�&m�n�m��c���rTD���fuk׎��q���]���5��i�ө�������XB�P.ET0r9\��ɩ��Kt�֥V�h�s>z˹�`m,�r�N�P9�n;��-C���(�{�huq�M�m���3Q9䨈
��C{)�rh/ETw�ET�"*��M������a|Sfu ��X�q|SFc���M�C4��7SCfI��>�IqoE�s�<��.�`�QB�x���Y��n�F�#�Hj0��yl�M~�t�޹�
ˡ�Q9��"*�3���7C\�����~�>ң!�n�v8�n�C�Q9�n�C�Q�H��m,�r�Q9\	���mETד2�;4�YǸ��Q�Y�Ƭ5�E
}���v�Gg
^�"*��@��W�kM�Yr�4���v���(Fpcי���2sTD���V}�G�M�9Ye�fP.�I�wE_����
˱�)�r�`���ڶqv�T̬���i�Lf�1��T�*+�r(�Eޛ�Đ^E*~n��Fu�4�aZơ@GET0XuTD幎��2����}������ӿ���ؗ/�������7)v{x�����i~�������z^��Ǘ��_��m���v]|�������;z�v�N5�4�>���>��<�s����x�y�J�'���~L�}����U�M�l�!�Ǯ���Ӵ~���0�bHf��N�0b�Yw��qL8�s�,8��=��FT�͛����C �S���;�$��v�5����)�Kw��:�ӱ�2f��F[��nG_nEf�&l�/�zU�	�������_:�|�K�ݗ�T�"�+bGS�2oَ�8��[��9��eǒ��i��oºd3NǄ��y1�a0�X�V��A^���kI�@)<Cʽտ� 
ʽ-R�	��fJ��h�y��{t�)��-�8P���n:ǁ�Iҝ��l?l9KY�؏�de[�>ޱ�S^]���r�;���Ǉ��pݸ����! f�u]d�-~��V�yr���Γwvo���<y��H�Γw,�����;�������̽�,��4XP�e~�O;1��)�8�&֣9�%ͮ��b<����-$'���w��/����B-S��,���C��Y���BXύ�%�3Z;�k�����"��<($w����Q��(f@��ɏOg���x�o��п���C�6b���������.(�1�o�����lp���{���}���{�[���?����������Wx����ݣ� 3����{ oU�38͌A�>���`_?;}���j���<I}�]� D��9��m���J��!�	|(�J�M�xt�u�Iu
�u�I�[� �<�����)v�2T���֏�IlH�w� u���(Y��( dw�(Y��O`Pq�Q@P�oS`Pp/U`Pp�V`Pp�X`P�oZ`P�/\l����.���/��з0�"�&�1���w2���W3��74�"�&5����5����6����˟���
��W�����ǽ��kA@ip� �o�W����Ͽ�?ޖ�}����m��W�\�)�w$��q+��y9��yG��yU��yc���/����q�d¼M�G��T�G��[��w������?������~����������?������7-� !P��?��d0(�ud��,��g.(X��ˮ��+��-��W��Kѝ�tG�߶���������d�����?���-���勸/�������>���e�z����>��^��'Ξ&u�|��kb�P�.�Ll��Œ��MB]�`2Q�I�K+e&
6	ui��D�&�.퓙(�$ԥ�4���4�f�`�P�V�Ll��ʚ���>�� �OC�[| J 'ʧq �(��Jwp�8 ���T7���8�Z	�[�4.ɺL<Ą��m�4"���ӈ8�U��� o˧q��ff��� �W�/��J��8 �W��|�� ��j�^�O#�� �ʧq �+��J��8� D> �^`3˧�RQ>�?5 z�q�d�^�=��;#�1Q��x[>�*��q ��x[>���m�4"���ӈ8 ޖO#�@�_���-�ƥ`�js�j�A��W����Z���ӸTx��cy���:���ӈ8 ΗO�r	;S�c��b�'�n1�BX�oc��c �� ��O�R�����`�˧q �/��Jv��O���-��J�~�82샂k��GvW�ڲ�,��z^%��H^F�Y���虺��p��;��R�ɾ�S�'1m7+��f����Y��@�f��� �`�`�a�_�Ȁ������#0��.X�y�����b6Y:�y�"�������g.^X�7� �l�����5����������#0�t���b�n����T���a:<��!6, 4BB#L�2D�*`��F�-�e��W�	�0�F���a:,��!:n#$4�t�-Ct�FHh��T>Z�����o�w`d�E��<�F>0m 榨�a�F�-`��F�nr�e�[�	�0�BA���a�A��!:l#$4�ۮ���0¼�-�etآ�a!��kVh��0BB#LW��2D�-`��Fx�-#Ct�F��a泌[���,���m`������&�gU�aK��V�Y}8]�D�ŀa�쉖!:�#$4�tQ-C�A1�I1tc�Q�AG1`��F�.�e��b�	�0]nF�ŀ�m�p��au����6 s%�j:�#$4�t-CtPFHh���>X�ŀa�<��!:l#$4�T5-Ct�FHW	
ϔ :���(&G�� �n��Zh��o�������j,:�#$4�TC-CtPFHh���	Z��O3`��F����e��br��%�y�8�A�Ԁa*���;�Do�w���i0W�ǡc0B�@�r����8t�FHh���Z�����SQ�����8ԡc�0� F���������ǡc��q�	�0C��a*���!:�#$4�T�-CtPFHh���X������S�<��Q!���h��0B:BX��~��JrY���Y����YY��n���Y����Y����Y����Y}���Y]�Z��
���Z qM���n���&�s��v��$�b�:p�q�6o�V붸f�7.�%�5ۼUX-���ݸj	p�g���� ��S� ��O�t�vSǡ��S��S���'ǡ�ro�9�6�q��V�"ϡǵ��O�&�k�yg�Z\ok�U�����:����lo�����͖8���V.�y�l�͕8��F/k9�(��qsy#�Z\�����^�(���7@q*����F��/j	pw�n�� �q�j	p��s�g���d��&{�%z�%�%�%�%�%�%�%v��k��k�!��2�n�T�,Jm�0�E��m�5ۖk�-�l[�ٶ�4-�l[����:Ўk��;�%vw�ĹT7/��:�X�Ʀ�S����'=oR?�{_�
I����񁪖E⳸��
G��ʿ��K��[m5���W�Jes\�>��D�w��� +����z-�Y���UM��X�R�E�^	�p��A��fq�w�J	��ի�C��l!�WB�1�jz��Y�ihVM��l7U/����� Zd�X�V��D�YpU/����� Zd�X�ܭ�D�Y�[/������ Z�HϷ<%�����8���vo�R�<;:~n�dY�z�`9>j�W��,OT������� ��Ƈ��Z���J�r�6NY�H��F��Nd y#0��=O��:�现�pYի�� F���QE7�z�]�F`.{&��% QT�հ� F��\���ލ't	�UtW�'��% E���	]�D]�	bt	H��<�eyB��\QE��z�]�E`.{j��% cT���� F�l.�z{��蒝��ZO�K@���a���d�*�~����eUs�z��	��OE��z��3	�����&�'t	��T�A�'��% �����	]"N
��
��
!�O��>�=��G�}��% �����	]�>�i�	bt�q��y>��VO�{�Oh��h�[O����]JI�Y �ǼӀ�QE��z�M�wQ���L�7>�Z@
��q=A�j7.�S��i�QX�&�����'T�Q�@35�N0�L�|BӀ|SE��z�Mo:⮔���i�Q���]t��o���������'t	H?U���'��% ���K�	]�O}��	bt	H?��<�~B���i�j�j�+j���Ku�T�=:�t�W��.7��T5S�'�Q- �T� F�y����	M�%��V���\M�L]�O�v#�ļ�f����	�L���	bT��`ꘚ@'��L����'4�N04�?��<���i�i9�ML�`2���L��%3ML�|�� �d��&��7�$4���Rm�l>!zt�ɢ�M|.	�%��TճO��o��|�KBsIh.�F!��G�,:����\�K�QS����u������ॐ�	&H0Yt�ɢL|.	�%��T��
\ѣ3J�Q�sIh.	ͥ������B���KBsIh.յ�W�蜑E��\�KBs���\��Gg�,:+���\�Kum���C�}:����\�Kumc�=:���y>����\��R'D���8tއ�%��$4�j���	ѣ�>���sIh.	ͥ�6V���q��KBsIh.յ�W��*��2؈:��B�輏�}:���y�����3`�	ʹ��v�j�r�4�KBsIh.�F_��G��:�6�}3���&4�j���	M��B��sIh.	ͥ�h>[/z��
ytV���#�
)�iB3�6���:I��I">����\���'D�Nyt�����55LM�sFL�u��f�}3�vh�^|��<5��qV���ɛ8Vο�.�h��n�E�LP��;�B���iZ[4�N�ڢ�wZ�Ϳӱ�h����e��6@��u�k	pm0��]K���~0���!	�6�غ��d��u�j+����avn���<F�6LM�m�~��_L��=�h����zQ�������47��\3O�%��Xw��E��<R�M4�MXB��Y��7�6n�ƹ]���{~��;�OW=F���^�U�Ʊ�M�,�x;��4���@��;�C��E���6ꯋV������=�ل{�/���v�"uͨ�X3�f��K���e��]����y��Ƅ��Fw���P|���#�g��0����;Ϗ��vݤ������Kߴ�lrzXLz��x��E�Ͽ��D:�1�z����Ͼ�tpMڠ���0�yt����4��;�ñ;ƪ���v������ָ.:뮧eL�Ԗ��܆�<��a��V� �߂�ag���yrjj�}�ui��!���9��܍�!{Cr��b�ˣ�m�k'C�eh�[BcEqW�6.ǣ	����*E��x���wL�h��}]��;ۺ��wvuE���E���E���E���e��6@�ދ-�pm�^lQF���Bכ�!���I����K�ŹiGkwoQ2����ϳ�[�ƍ�����`�������-������m�ܝ���\�r͎�-"��~vgA("��~vg�{Gԛ!�/�čL�{	�T7��\;l���ld��媰;�"r�*��F��܆*v쮈\��=3."����3�"rym�=�+"��d�]~�a�%+"���;�A�o�;�ˬc�ۨ�,qך�҆>zl�;��3�=�[4���-�g��Z�w�\3��m�b�c����uf���L��Ϳ�T}�G�M��Ye�fP.�[�wE���ɀ����ߑ_��;[��w���m�]�|3�#k3�t~4�M�Ϳ����M�=b��|?7m�S��v��0-�`6V	��J��W	��J���B��K��嫄3/����2�����"�/~�Ӌ�GT�u��������5����JT�4����}��or��1%g�$��N+ZZ7��O��20��T�4���K��KŷKm�K�K��K�K�KR�h��#.Y�K�	�/a�%~�Ĥ�8�\�&�0i�I3.k�e�x���qq��zq����e��,˗�Ԧ6�pi�K3\��Ҍ��\����f�4å>��i�O3|����S����f�4#�!�iFH3B�Ҍpm�Ҍ�f�iF�f�iF�f�iF�f�iF{�F�Ѧ]�ѥ]�ѥ]�ѹ?&�?��W������g�o&���o&���o&�$�o&�d�o&���o&��to&�$Qo�'��s[I�$ƶ�,Y@A�)�Z�ͺ$��`iW"%��{�=1�0��l�29��n/�pl�P�N��I%��Ɠ�R��B��?��!���������x;�`�r���戈�h'\+C�7i&"��!r��NXV��n 
7��ޙ�ٶq�S��>�Ӵ~�o�0�bH�u�>��ձ,����g�O=�
���G�Z�z�5kW'�3|�u�����w��nc��U�+a�"�|%4애5��e�]]d�5��,W��vq�o��"�9��]�4�z�/O��-ý�C����oݸ��?��ny��E���)B�n �]������*����2��殟�[��=����n���;�[�U}���э�64��GK�޼XQ��r���/C��ʑ�s;�
�l�dw��О�n��a!��m�t�Ո6<�n9hv�액��u�����Ks�^t:�8�v�nז�#:N��6")��W-N��!j���L!"N���D�1Q"��y����~��	6v�f?_�h7�,������^�S59�=�^x<�s&'����q��d`�3/<��9^����݅�8��r0{����D�e�x$��k/=��Bw�e�{������Ɗg�v�h6V;��+/<�Ȉ��޸=/]x��f��g`
w��̖��'`
s˻�3J�8���)�z��`�%��L!"��L�d�ݔ�]�*���Wѽ-A��5���"*����C�����RSx,��Jno�)<�w�ܗS�����7�p���I��>�E��z�����O:��<�d���O!��?����ǟ��'zO9z��>�OO)y�ls���P�~���=��r�O¢\Z�4�6�=Ʉr�Г()�%=	�6$�=��e��'i�\��I�:���l9�I�:��~���ũ��s��'��\.�I.:��~���墟�s��'��\.�I.&��y����b>�%�\̓\L.�$���<���r1Or1�\̓\L.�$���>���r�Or��\�\l.�$���~~�r��'��\.�I.6��}����b��bs��'��\.�I..��{�������6����6�$2���=���"s�=�K���7q���3z�vy������iE+Z�|ܘ<���O�CCƼz�(�{�.����>����T�W�;���F?�K��x��q��w��t��O�����w?��?��/������G�-DE~�����t��m�����ח/���)���\�l����Q/�����w�����a��|������������������������#�h(��~Z������{ �{�������w $J܄����]��o}�nD�_�گEʹQ�	��ǩ/���~v�Q��i�TӇY7Ɛ�gi��'x������x�Sta��w�_G��WD/mc|�~|3?����Km[������m4+������fc u��)��?L�0�� O9U��=ֵ� �s��=���� �|�z6�Y��>������&>�����n��&�{��oY��$CG�o⿽�X�M?���C��*�=c���?����Y&��1̵O�vXs0@Q�
�;���#
�9�G3kZ����_�vc�[#��Hk�ûyc�~w{�����y^_���`�ٛxīq�!�[.�'���-��/n�f����lC>���nz�S|��ہ�S|��ہf��٢h����v�����`�6~�%l�~K�;@������#�������`��[&�'���-�ﳰ��- ���o	�6~�%� ��=�D�����G��(��]$�/�zx46�mp�m���q�F�7�qW��3?n�xZ:�o؂��폗-��~��7?M�������uH�蕊�wo��w�RA�v��������-|{��W!<��.j��뇏ʈ���6�l�g;�m�H�ܴ��M��ڨ��]X5^"��m~����6��O�&�ܮk�M��&tL�P�0RB������h�7��@��R�T:Д>Zlo�Lzg\�e�\!=[HOң2z�������_�vg\�D<H[�Ľ������Ƅ��o�u~��]|A���ut4�}�����H��+�K��M-�z
�&j���f&��o�fY���4z}�Nq�s�n��t2��]v�[����2���ep���_������6�(�К�Ƿ�l�#�����M4��(�qw�����vM�٥��64�L��a���6���E�bh8�'SY����{i{�k#��+۶Z+K1�n۫�ظ�t�Xjm�>1��_t�Y��߄����5��uC��8����G���]#���]�_���8��m&ʚ��F�v��1�A���������Y��!̆��u�oc�fl�Tjř�N��K}��)��Rf4!��6�� 2��1x}��ڦw���?��٠�J��������ߕ��*֪��|=�����+�eTD���Q@VŝX:s�������h"����~��e�r�5���$��*����+��q������_��T�5}1�0������?��_���_�o�w��>CyҾt/}��׮07u6ݬ�A�=���p�{�(;�&��K����0����V]T4��z�К|g�1,\�-<����jl���xQ��S�����þ��_��o,�h/*�vvw�i����6��k�����<�ڲ�q�f�)n�У��K��g�E׿y�ũg���,j�5!%��!�?
����Z{�JEFuf�q�M�}�̤������lÒ�**��V�dnU7��_�T�B`�Y��W���O\�>}wz�
�����t�I��rs����#��������o�Oi���S��Z��z�\��[;Z��L��h5K��ah�oO=�����TNQ�ς�Q�/%��������{��&���� �b
��ꜵ�K�R�+(�r��E�u&�����Y�4mh��/g��t�+()pZ ��*���۸�����-��^��3��'��ʩ����c^~�L0����D&�$M���5���8���}yN�=}�i�!}�;{Cʾ
�����C���H����!��ځTc�qjz3�M��	n�����v���Z�e��z�檊�g�g��
�Ӟ,�$�u]w�����7��������7�������G�7��v������>Gk?�)�F۱oB�a;�45c��]����}NQ��}N\Now���D��>'���q�^�ׅ�qɟ����t�M�g���.�^6������-�m���ָ-�m}��ָ-�m���ָ�}���~_¾�*�=���Q��\F����^ތ��Ng��ʾ�S��-x�N�m�v�qli^�e4j�v�%��˜�����1��Vi��8q3j/��̨�O���x_R��U�O=m�n�M�oc$��%��&?7��+����M����;YQ	��=g�Wۙh����я�/�\o������/�v���ٜ�\Z�|>�ʣ�&��t�y�Oݸ��U���ĩi[��;�f;/f-ꢂ�%���C��Y6[���K�7�.Vӹ՝����)�κC��>�G�~#�KG޿d��O?�e�yRDk}�m��t�Ǽ�ّ��	g�=E=�|�J7���F^/-������E�W������K�����z���4�_K{��V�:�y��$E[�M�׫I�b��,�-����?��[��p�ѿ��_��g��������o?_&�t�݊~:q�O)�����xظ��ɧ��!n�1q;NѮ�ZBp�2t]vM������p{�F���v)n�(~w�=�X��lm>nܼo���E��h@�y|K�5p:��l�MV7���X�/]v��]����ͱ�E�t��u�}ܚ������ζ���@E}��r��]�|^w�O�u��?���Kŏ��\���d��~J�\��Fw1\��^4�U���Km�?��>��20��}���ϯ���i(]ή��-ů������s�6�~�~���Ư��?�ǿ����?��_^�?�.j�ͻ��{���^��e\=�����ŵ���ׯ���t�����Bp~;m��n�u�����o�5>M��r������ӻ�o?������?��w�{�ʝ������o.{��o�m�w�����|�A�gad�rk�����y��"��a_n�>��Ͽ{��he_�`Z��xA�i�����"�Y3��
�}�Z�4�+�W@�qr��`�)��e�f����;��=��@�����cOL(3���0��2K(V�ab���5n�;��mTydK��A_i\�3���̦=���z�i�9�ٳ�V�4���;�9Tn(���J:L�\�m�6���r��6�_���;vI
@CY��[�����^m(e���|Xoq�E/�-�P�;�r�s��qtG�q��~�իM�,X���n3��r93.�W4!}���v�0r���9��FC�~b=��T	�<ή7(eÞUi|>,�?���m������}�&t�>y�z�>Y�\�v�t~\�>�`��m�5��P�٦�2��Ն���//y�l;$`���Ѝ����f�[�-��k]w�Qy��{��di�5��¬� ��l��6�����q����gA�n���Y?Ka�W�)�'Ǖz���^X^�~QЇA�9���P�����ϑ֭m�hس���^H����e�mpj��ur�e74��Vgxʼ�j���j��U�ϵ�o���*�5���^�VU��]�}΁��+]���ǧmK(��e,x@�
�2�Z����
�'뗽�u��6�]�þ�]!��ZЮ�if}Ʈ��j�1���s�l�n(�#x��L��"x#�m�����]��Q�4v7�±��R�n�3��`E��ԨҨ}���-w�䋗.)��x��:=���:&J���ܙ��i�����xس�r���9vzM��Խ�����m�zt
+���6�Z+�����#�^�*em�v��N���
��-���a*�>'��Q�/�.)v��u�OaE�������Ke�\ߧF�8�"A�ۊ��r�Q�SX�F�?�T�=S��䍺ף�M�X}�,U�O�Vqǎ4��:�ݝ��ҩl��2����%<o���Q�n>�q�þ�ľ����þ��۫�*��<�)l0:u��T�ó2��j����X'r�Y�}�nmC�0�VR<��ލ��5A�%\Na.a[p�_�w�,�ǉly�č��ur�[�h[p�MCmgO�+��.��݄4��m:��p
l�9w��-{�Wô�\-�ե��a�*]���]}�·m[�]|?��	��c����UG����/�	��<��ͺ�?'��'������M��W�kh�r5��
�˘�dIK��ע͏I�=�[��+뵕3z�DfW��
�YT~�,S�Cf9�����s���kͳ+3�s�J�z�8*��éӤ�8��*�:M��究U����I����af�HXX�-V�*������V)9������Z�tE���{}��v������aaI���û��x�
t�G�W+�ڹ�[:�R�ָm����39E�-;�S$ڊ#9�P�?u"�Y�	w_��q;7y3�����ž�eيD[��J�>@<k+r����vs��+�t\W���v ����[�TP��@��I��]��@V�h��R��|ܶ�{�,�F*��w�ho)���R��kI��3���έ�L񅅊��(ɣ�w�w�bT�W���� W�(l����D�'I��g��j��
4��x�*?9�� �����Jq#A~:�V���w�Uk���­�ᗎ�a�ӏ[��-�?�d��]�ހwH��g�S�`�v�COno{5��Q$�=No�v���G�0��F���[�ހu�MET�vg�\��[�>�V���8�S��KPeü/�ݔ�Z��Zd*�2�`�v.1����x��Q<�=N��r �/��|[t�;���?�k?a�Q��(Fqn?��״���ö����e�������|�W<!q�ŉ���+���G���Y�*ܶ�91��lĲ��Fx�О��^����'?J�Ͽl������dYY�a�ݮɇ}E�C�\f"���O|�@�6����-��o��V4�}�Ou3+ŉvC�>��+�)9�D��\Z�R.���en(Ț�tB�^�Rg/�T@���>C��Tț���q;u�wX�=�H+Ȋ7*��WUƀήY�m;���"ǒ�۩4���C�V���D=����ڋ�׆Q<n��mf@"e2����H*���H<���Ʋ^����5d<��u5��0���7���c�q~�����ɦ>\����3O�ؿ�Կ��?����c?��ş�PK   ���T7�I� �" /   images/39ed726b-0701-4a7a-8bd7-442054548109.png�eT���.ڸܥ��]�C���ָ�&hpk��-�-��$��`!�Yk��������c�1�=���9�y�U5߷�yXz��R����� V���	 [���� �  �ǮM�[OOWAvvg6s+������+;';@X������	����9�P���Y�P��*s(�JBl����!��*Z���V�b��¾��N�NOs�������������w�S�0�t��V ��Հ�.� �%7����������������񜝛���_��K����E
�[YjH����%B���|||�|��\�m�9�9�ع�X-X=��=�}Y�=h~C��!�t�s��sq�n�[�xy�PS��f����خ^� [Y�C!NgO�Ǽq����c�v6����ߦ�����t�u�t�uq��G�S���(��i����;������zxZ�������'�?ԅXhz�{��?��ORA������������t=�g(le)�g,4�L+����֟MG�ߎ
:�;ۈP��ZA�ͽ=�E���D��O���+�0�_��흥;�����_�ӄ��ս�W��w������&���t������o���x��{δ=�m Zw��y��ӿ���U$(�g��.����S�������؁�ܥ}=ͭ��kS�]/i�����u���o�j�.V������ׂ8꺸;�������I���_�?��g�����R��(S����%��Y�C�������?$�!����HP��!��x��y<B=���8�z�j0p |x8DT @) x)  �0�I��p �oy|E@Bx|� "  ��"#� #�b��=
*::���g��Ϟ�S`QQPq10p	�1�	�����������ņ�Æy�yt � ���O���C@D�G����E���  �6A�����W?6"P�
�Ì��@����L�u�������m������@��M 6<'X�h���f���C��O�JÍ��aZ��!�~F2��y�wK���,ت) ��/�aS��\�
_���� `հ����yTs���́nj!�Eo8��M���o�>� ���ņ�~4;)�[&�{ݟrY6���d�?���F�,F�r��X9n�T��\��R�T���'`br_ø�G�6�\-<�[�;��8��/9�Y)�#H�����Q��J���N%D��f�
���Vvkhh��M[-�t|�_��Ȋ�/���Ohy��l�\z����|����a�6\i�7�?�(�7�,T�~�=�<<_w�=Y�\Qu���fV���Z�*�tJ��ѝz4�e�ut�k����Fz�-��F�r��EV�����e%����?�Ԉ\��z�v���c#�~q����.�#�*�M�1Gy�z�.�O�u�g|�H�����L�,�����>�����V��ѝY��]'d�[�~� ���w��p�y�3#Z�~��im�[��;�r���z[��ر��Q����5Sc�C��iFaN�_g�5�2���.��Ύ��+�8��n���z� pR8��=��&C�ڽ��2��s��c_g����E+�� �?-�
���N���p�1�������P�{Lc�R�em�������9kb"G+{^I�{���n]כJ��J���Y��X)"@��a�A8P��Vm;/������=^������=���	��/���dW���������T f��DlѺ�R�n���W ,�Ђ�b��6whug�fT*Έ�� ��q�s)e��zb�O���1��̄�R��w�M��&W/���Ų/
'�=wl��"�@E ��y������3{<�`E��45��O!�� �����%���.�5w%�?�NǊbޟ�Ei�.���i�{�ww��|�2|���~ T���s��`N���!L���=�}i�=RH��h���eD���GU����W"�G����|�p<����$?&�|6�����m���	�Ӽ�c��jHL�e}>~^��b��pd��b),2
E"s�l�d=�_�i��}f9!���)�䳗&CדHk��zzv����2����u0ǆ/�I�	����`)����l_� [��X\n��0�dn)�����/�r�}�@��ZY�X)Za�'���N�A��` ��m�
z�������$$(�N�PE�cJX>�;��<mX��*\rz�N�Q�@�h�d�Z\�U�(�������h��c�{�Lb�@N����m����o�x�����@zw H��| 
]�3a�s��/�2c�K3P��>?��#.̤e�d_t3Lk��P]����}��:)	O�5ɸZ� B#�B�Gl�i���+��D�h�}�Z� $�㭛�1��M���{��;*)P%,j�tZj(����:��D\��<�Px��S�9��]z�Q�:N'oD �)J��3�r5��J��<-��`u:�)y��3���'pꃟW�q`��fUB�'���J��5�c�P�.�I�~�o����)���:Z��s+�.������S-���K�.6�.k���F�I~Σ^�7Ŧ��8��j��ĳ��!��`�" ~Ҩq��Z �*�-h`T^w��v�#��*&7��j*�1����Z��[���24�uMEִ,K0�iALlc�ٵO�HȘ�*߾o�ߪ3����a�d�O����u�E��H�I� �l�;�o�g��"V�ܸn	�m_;
��AVN�? ��hF'G�����M�Y���r��G|̌�Қp��X>��,)����tG�]S���>�����sK�seA���V�bZ�W�s@��4�����۹'��2���#�55����f���8l�)���w�m��oPSx�/��R3r�4`JY�@b�p�)���F�׺lű|��<�Hؐ�h��b�Q�H�ܓ0x�}^�9�/�1�&$>�����w^��'�b{�}��6�/Q�=0��ya�5i�(�����5K>ׇ��������t��7�b����������/���!ž��N~�v�'	E���ю���R�od�6y��<g�F�����:8��;Yǵ��8�Ѷ6f��a�d2�]���9�&;xaJr��� `=�I+s�c��v��m��e�h�79�b�8,p�*b�W�1� �4?�=���\�it�����v�pt��"��y��u�t�|��Z���V&�n]��.�^Nt��	)�vu�~�[�?�7��y��n��gb�E�?��|���îpg���6n>�P����\��b�q~�z��Ӑ1QZ{���L�P������w-+-����Nd�z��f8]qpf��A��J��8�4�Xئ��A��!H�.G�ÐU��.hmG דܺ�zo�ɂ�}�$��6	r�`K��<p�p]��[7��;���꺑�Z�e�#p��ҍ"��י��ϴe�^e3�[a���*0 ����ZA!����o�Ȳ��2FQ��u�i�+�jA��Ղ�~+�9�p���A��̎��%�y�O1q[b��X���A����
!g"�|��� h(JL�"��ړ��d�*�٥��a��X�Q�@ 
��2L+�i0�7U9��0��{�����P��f@:�J��9 ��,�A$��搘C.I���+k�Ǯ:��H �v�� �6��2�h���2Nhh�n��e/0�]R){f�>���F*�j���������o�eϧp���՝J����[�����I����{�5�'��s3{'��)E�5���³SSS��l��~e̦X~���C��y�4�1�Ca��66{����Wڻ�����KF\v���r�C�K�'�C>f,ot�}����s�GKw�}�l�bŪ�����) ̾���<��45�2�Qp_�4Pnq�%=k�R��X��4eט�:���pL{�{y��㵎��$��==����@��r���S��E9��{>��$<'�Ϋ�9�9*lE�$�J'2��;�T��Ur�f;z���D�K�����k>7��t��Mѓ��9�kS��oo�r�7:�\�s�]=^
�*��s�伡�v�q�A�#h/�,��M�Y��k�T�u���J ���^��������[A�i����ɻg�e{��%�~$���\OCA,�@��j�S�O(��mT3�M��VoVc��@]�]�~�=�w��Ӵ�b��=�Jq�����+k����Ȋ�ja�+��耙7�闧&��)��I�#]��	�!�Ohto�sP�2���m�����(E.�?ʁ�Z���\����Hy�
��y��q�͖@�w�[2]�G��nu��e���ނð���<"�_���ĭ�"w�g�P۔8\��zO�<dd`�-���t�g�:���Am�l:�Hw#�����8p'+��(4����w�ߐ+s^�פ�]����hY����ۂb#�z�V@TA��_u�oF��������bd,�(iX�d������f3VOm�y8����j�:���q����
�ޛ0��؇,
Z�^e�#�G�  �+�y����Gq�e�e�}ty��eCm��6h�K�?@��9&eG��%!dpy��=��8 ZB �~X�KEEf\�nϠ�n�O�?E���>���!�0�y�J0���%`b��`�C����H�z$���)�8Wއ�gfh�\zM�'�aWۃո�k��Sqnk��``�J��:N8������A�<h'�9zt����h��8�$�T�ڛ�ŵ�ST�7�����Y��y�uuZ��`��ҳѧh$�db��'�9C�3�#�ll�lc2��)}�Y���Nb��x��s�6?K2�������@]�/xz�-�̄Q_DGׄ��r"�Hw�n��',���wZG'�����mY�Z��9+�q�^�厜[�;zM{--�ݚ������m��os���:ږk��W�$Xj�ղ@#3s�c_b���sԔ�˿����4��s�� �y&lH�`ۜ�2���]*���o��`�w4��S�~B�� ĒX炌�@>x3
����b/r6�#��L�3a�w��e�2�ec�-��nw�o&k�'�:���l|���Q|i`�Ͱ���\at��,x,Z�d9-�e>M��X&.�썧��Ą�yi+0��c�Kbp�2���2kݦ�Pgwj�W�35·���]�nmz9D35�X3�V>�i���[�F(��r�6�E�Em��cm?�_pF���bfF@�9>�k��ˬ-/|�'�噊� ~� �;V^Pi�}X����Q�T|β�N�N���[��޿�>#Y�>Z�8 ���"T����z��c����h�@�2����"e�� �iAPX(��־�_ |-��3j���ϵX�j�l�?�^12����}F4F���U0 O��Y��2����8��˥7���tCƿ ��3c���)���y�ð�1"��D��-�F� ��� ��ŐW7���ԩ�G�TӶ;���]8�h*W�A@��@�P��0�B��S��ꇱw?��'��F ����8���������p^@ǩ�d"|(��1���QXx8�rԅ���lVc.O��4�`�k�]}����I�+����9���O �9�x����Јe6�xx��ө����g�l�o9�K:&P���9�nz�Q@�����+v$@U��@<.�H�=�r�F^,}�4'έ�ε�#�&�<�1��`�_eT7`���{tEN�>E�>���1���Y�85У�#�π������d�u2�9]4����Z�6�������f�aۿ캦�>j8��#�ݺ�Pa����������I3���UHV�z��X[Zn���y!�����m�q�_���j�7s���9��.��Nm�����9��������`��֞�gL?�>��H��Kg�Ծ3�)�t�7e̯M/��3<�ڎ��~n��M�ٺe_dE�TG�N�UR���;f�z�(Trs߸�ɜ���{���ۅ�ӎo�O�)[5���d��wV�j��:�����J��J���o ZB������\ɥ$�)g�l����ɤϰ���7�;3B#������3�w�����Q2�.6��YzC���B��`c�&�_�<0щy��J�٦x�p�<g�g�4�o.;;�(y��|�?5쯲�ԮzxU_�Ld/�Sd����i�CѬR��RS��L�2�O�%2+�?��p'�P��~ �s}k�>3��!d3���+r�ڬ�n*'#�ꆧ�`����Ƥ�We�Sh��Wo��V����V�q��ĩ�f6�G~��GS����Ю���<�_�b��Ϡ�Ȇ�.d--C��_�l�Q� 9������[�Bl�ZƓ�=bW����6���}���1�'�ּ��ޢ"�.ES��"^�>YAΤT5D%ӆl��.����
�hV ���`y�8��|�Q���k'Lx�+f�s��DN�ׁٌ.*�;�qW"��?�<([��􎆥��qq!�Ux����8�B)�}v��ʹ��o��G�@����U��}��Ϣ�4H�0�K6�r�iE{t��}K��ғϳ�_[j`/��D064A��U~E��o\��40֐'�o�����-k�l9���K�+��-�&�T)�
��w /'��-GC� �FS}'`{s�`[]qxg[ص�����A�n��W`t�<�Py�b��S�w�����������:ZZFL@覱��<�k�6^�c�V�a�0�{��A�
��8��i0�4
������ U ��]�B����y��@��� 왴b*� `4f�[50)�du�1�����{�y|�~��/7��F6r���e�����BOP ^�=F��֘v�H�������X
xu"2�M��9��\��􏮘#�^�]��������|
%G�u�.g�t_,�Ϯ����+�*���|��Y�(v;ݍ��%g
�b�k���������H�t�11s��Y��j:������[e�o�2����M���1BF{���������s��%6#� mn��oY1�Ϝ�Y�=r"(��;4��4���V	x�����>�:\�
R?��-���M�T1KTpbh�g���*��F��(�uSCF<ͤb���[ap����8�i��u<W9q��e��շ,f��X�3�^T�\O��Ym�:u��p�\���\I	�o�����ke�`f�z�_O7�>�|I=$KL��gё�Y��Ě~�Z���M�kZK�I�%[�$��a�hG��N�MղO�â�t[�v<�L��*΍�Q�ĥ7��N�����p-l1&n�`��T�K�o����%x���Ƨ-+p:$��_T�Ҍ��$7^��#7> ��,�q�������
7�[{BU��6�����3�������	1t��E�*���9��b�џ�vB�a������s���p+T�#�i��Ԅ$�����z�{��z�����KQ���Ur����,�R�h*�$S��3��y�o���
/�,�7L"���-⭮M������,��Ue9���z����Ɔ�,�եq^"�(�o!U��//����١rw�S�%��N��<>�l:�O�X�@��Pϲ�s�ҫ\p�E�^�8�kH��{�Ȳ��8k����Z{��~}���Hp=���b���t�Q�혬Lg�P!ƋF�����1�SN++G��[\�%!�W�m�c���	�����E�j��CGdט��"��j��^��
���	�xF_�x����|]�����<}�Urr�#��eӌ=6�Q�6��3�8�̪��H
Evó��9:6�.��ѳ�� ���J躕��K	s3�R���Q?)W=�YҼ)�Bi��iڕ���[��KRGe�k���K4���u��Aۺ�C*�����ab%�2�|�����Q�j��#�_��g�h�өJ;���`l|rj_yh�(W**p���X42��۞i�-v�N�k+VEg]�2NO�/u�h�����p	R3ʰ3�q{�gJ�F͇��v���<�"��2�����Ѽ�-���ˢV����#97p�j�޾�n�(<�p�5�n�G��D3��e^��Hb��M�ܐ��;L箶����}L��b�����hI��3�{+�������\o�Ǚ��/N���h�WoสǄ.5��ӆ"f�S���w[��X��P��k�_7&����|�SJtH�=���SV*���� m4���$+�m��S���﷜r#�r^��*gF:k��s��溜���qBՑ���>���0�b�H��$#g�蔗⫹���}�alIa&��2�5�T9�R�n��
�k��3�옘��2Y2��J�1�<���n$��[8����e�/��?����_�ھ:>��l�cM������CVlz�@v_׳#���G"GEմ,�:��l����.��*!|�f��Td�Up�թ�(2x6FC�D㖜q������܉Gl�r_Y�����> ̻xQ &��<I��S�1kV
Q�Rr�q�l��l�j޺�4Aj_�^�֪��^��`��U��ID��#&�wI���oa�x�1��Q��0���J�g_��V���	7j�<i�+}�+�"~n�.�!�\�3I�[�pBR��o{��5����;��Fi}sz�iu�d�\����eι�L- ���Ǎ��n�-i�Z7�ZU�	Ym<_4��EG��Um	�k��푆.4�^��Z9���x�t)���`��U������6*�m�97��A�4��ѺR��	��,۩�1��ɍ����UU�V��f*�c���lӧX�p\>sN�&�Y"&S��b(i���?��%�L5�~#��|CJ&�w8M܅���@����.�N���.�5�E��u����'$�Υ9[oj�֫|�ݷ�ry�G�`Q���w���ˊ�҇	�i����
�?->���`y�X��:�<W2j�N}�U�R�Pߥr*OC�/�vU�P��'�Z��s*��{�7���~<�i�:Ѣ��_�����@m�eAB�fQ�*g�BՍ��W[��'$����8`��w.>�D_�RTsS%T3Y$s���:�I���ܐ�k�Ys��v,�B�T��B617�R�ߌ{���A,!�Q����C���Z��c�,�ZbվZ�98�����_C�įv��*Em}����u���E�m�ߧ�ȓ�*��|�'�.&����jK�+�|�hM1�Z������-I&��֏m���<BŨ��
�_5h�q��t�6�D8��8�U��? .�QLM��;���͡3|oVL�5���s����v���G+I��/m�QI�W���*�K���(�sɽj���]b�-�^P������� ߨs���t�� q�xS,��ѹSLh��\�}i�jχ��IU���si~����u�l?�rG�j�:pჂ(eq;���<%.����3�E�`�+�$�����\[��-�vſf�Fɛ�,��gs����d�ؤ6c����h8�[�
��96d#?�[�9#�EcI/�,��USU�h��WJ�4���;�� �u'�۔��fb�BU���s�cNA�xcAm��ڑ�qU&�G�c]���/�
�q���uH3��y(�\&:���Ӷ��v%t;J���.L�'�sKe.�2���o��KH����~^÷�H�:��Ag
<D�MJ'\���g���+�ߖ������~����c�6X�?&�jk1���l��E�al�}���=hO�}=�Uz��ޥU�7'�?+�w|ݫ��*Ѧ�$ZQ�"�Y�Y`o<�u����k�E��I���zu>Bу���EL>�수�?�MJ���b��S8�ތ�� �K��;�[X<cc3._p�8K�2��rkx����"g���O���Z�I�T�c���+�<��?���kW��j�4��= p��y����z���:����8%����BH��cpVI��^��GI��,L�r`��r���M{�z/���}��njt8>O ���Y�h�p�ƍ��"�'C���4�\Ǆ����U?���m�B�Ա��FmJi`\���,W��жqs$��0��;_f��G�0�ek%���0=8�C�{Ԓ�������;��a�a�_�7VB�c�$#^��do�)��L*B����=@a^UP؄H�h�~��(�w��	%���L�=���q���E�,���2Eؘ_���6�縮F�A'�	sRh͛��a��~siR�5^�$��W�f]R].�?�c1uP8��ݸ�5� I����Yֵ��
O1�v�Av��3������6j\c���J~߶N+n$����6�>͘�>��i�7>rJȑ�Z�p@��'��E�M�}�N��׍�(��4 !+��'��J8���:9���� K
!��I�g�W��t�_P�Y�+2�UW�c�F'/�mγV>���Pܟ���L�A&��g�s�G�&����jT�MS��
o��ջ���ӦV�U{�B���|V�s '^Xק�tݍ��>B�sf6PC@��	ٍ����j�K�]��+��r�/�_ pz���+�D�f
���zv��
�#2�n��Ջ�hܪ�vgJ]�1cj��5���s��.\��99�Y:�kG��-�L�`%}ȋn�j�/V�$��K*V��pM���d�4��>o��-^� ��H��8���-���@պ:뚅=�#�p�.}&n�ŦKK�˪./l�no�	�3>� ��.vQ�ׇfv\�FbY�L\��;��y�>Q�6`gک�6J�[ν�����	E�J�wkwxNC^�Wt#��Gv��1j$��A��3�p����Gp�Ki�'=T�[�q+��T,~C�ԋ޶rŬbX׈�;.�E,�0�!`j.B�pX8�u��O�_]�i���X�?"�^͎|-���=bP/!���:�Ҩ~H(L�u���t�� ������jEY!ɱ�,3GH;���T�RDҍ���M����@�6�
~KN����`j�-g ��VL&���9��uc��Y�ԫ��h��u�t��L��Z�n0��W��Kp:E�1�c3�5ŋ�fƖM�.��H^�"������������EX���Q�W�$C�Aɾ!TϑF���XL�C��IH6+'rX��� ͊P{���p�ں�J��v_�S&<R�S KliB�x�"�ey�w�Z?�8*�q���d}k�ݎc��<�д߯U��e=�/Ke8a���tya��c���b��`�k�R��/D�W�&I�m^5Fʳxz �rxrGJ��?J;��Dn���_�5U��7}��3��%��9�,&5�mAA��/<ێw뫕	黾�tt�S��Z_tz�f���<�~�μKv��929n'�QjO�4�8��L��|����Z5_n�K��x~h�ԸC��G���+s��80��>��o����2��;�S@����kf�%g��KK���䫕*�s<�ݒ))�]N��<o��ێ*"U�)��*��g��<��X���;��3��AFL� z�OX�#�t*��3u�u`�Ɩ�AԮ,� Do��n'JE��)Y4\2��"D:�P�g�u�3��b��2M1.'�:A1���9��N�s ����c�7���]�g(T���Q�x���@(���T�6�R4F@���-���p��3�)�/��|�d��%�9�VYu�8�Z�2�K;H�ԃ��ͥ��ڏ��壪2��F=:�It��0��u>L��}���X~�M����'�"�9\w����d�<ؾ� �e�%��P�n��"o5\M���gHXZ�-�Hy���J��T���Q��kX,�U�k$w�.Wꉱ#4��.[�Ѧ	F/��.ҭ����o��m�L��� �F���+�ɯ"�Q��w�91�pV��"Pq���3v@�;2��T#Ⴞ2�z�).rc��蠢�Nx�椸c���kڄ�];�!�1A�p�mP;����|�@:+<+� ���-~wdȆE��B���`���ʷ�b��pp3,����Dp�W��T�R�c�%`�d�2�p�:ud%qۚ�6���� ���8����?Zf�a�E���n�;������嫕�es+1k4r�ӋR%������Y��ߴ8~�W���˖.^�%f�YUu�*�*OZ�F����y7Z���C�Y�������rg��XKB���.�>o�J��.��S�k*����u��m�C2��pG#p��j�} ���2N�d�gn|[�T*F�2Xx���owM�_Ӗ8��j⮓ߝ'�V��>�"bo��a~����E����,��d��,P6��H6��DH0���a8�k)+�>S���6�2�M�D���AE�ĻͿ�޸K��
�q��i�q���� ��x���_��U/>~	�ţlU��������33�o��˲�lX��|?#���U᭏u��A%�uv,S���ʻ�ϋWf���;3�b�2��F�7�;����	ϭ�E	^�'�}[�#��DAP�ݞ�I3*)�z�	�u�8n���C��zcf.j����)��C [���r5]q�����q�KtB�'č�4*!�G/�{OL,qU��2�ը�a#x�(/eg�}F����)m�H��n���m��߾:,R�����|	Ѥ�������,#ۡ��UO�z�^d�~����^o=�e��cd=ia �b]�J�m	Jt��o��GCyO��Y��!'NA�"*�WD��nd�"����.d�E������K~��Ç�:�y�Q� �^���2���h���j������W~~��2��I�9��{)��og�F����202=�/k�v/���U6�,3�Ha�RH��T� �����B�[�&�T/�Vd��2d*G�A5!~DD5�$u8��R�CN��KG�F~����
����`�,UJc%���K9I梙r���>��G�2�H?�Q�4�9|�9�ZN0�uG�G�^��Y.��y��@J./��M%~3��6+
	��E��)�-�s����<w�7@�=wP/�GE�fq�0��8�J4T�J��b���uҎ��} �Ҥ�v;}�e``�d�+c(�||>�`�i����{��0�P����s��������b�2���;��D��&��ʼ �9��t�_��1���RT ���e��qR�Z�_'�aߏ����ˣf C%�,�b�WJ`H`��j���	�#�;d�"隨d���f��
ѵ\�\Qf$k����!��׶"L��6B-}?�+Y}�2�"5���/9��	
'�����Q��x��,�&�Z+],O���S�v�NoD n��.Dx/[�
a	�yq�k��[*Oy?���][�i�+v�7�V}yXl�W�N�u2�:}y������9�.6�ƜE���W���Pj �1-��ޱ�k#���<msk7��j�l��h��';�{9�8�����2�#���=��Qq]�w&��������ܒ�5%iu!o?t5=�4b���Q�nX��X�����Ȫ�*kf�j� ~,�-�x숝�~���.G9z�36�Q7��6��#�U,Y�I늺o�Ky�ʢ��'qҎ4�)t��r[T��L���݋
� �ghГ���.���-�Cݜb	^@�hu�c���q�X�L�4��4Y�4�lS/FN,H��9My�W�r���Iy;R��~j�@�֞Lf��Y�vpX��� ��1�n��0�h%������1ᛪY.Q�[\�f���85�m�Qo�h�γ[
���=��4�܌?�nc�l�T��C��▖��[�؜`/w߾k�j<N^�ަ��ϱW�B������6����ZH�$#URW	Y� $4�0!����R�E;{�J�
�}���b�\s~�rP�+��o%p+��3��v冚�y�Z5P�2��Ǫ��i���Z����+R�+E�+�� ��[fHwd�8�K��+��(#\,�;�+$�$e.�Z�f�e!�
>�/;�v����R&�v-7|���Z�$�$�??>�0as$�z��h����~�Eh��m[������x|��L���~;�Q)J.��mr$�Kf�Tuz���c�D?@EV9�&,�����O�V�b�����P�a����Qs䢲�"%��8�f��ek�L���fI�f�^@�{s�ڌp�]�]����6g��бTC��4!2؛kvf˺��'`
��=dQ&QQrhh�P<U�g�l���wJO�>~�07
�g�%�9����r�z�}�����7>%�:���Y�����.�������	n�n�v�	�v��	v�v��!�aْ�����7U$�J�p#�/�߷ڪ�Z�,��S�����|;���	����+�0nxf*�Qa�C�F���47D�	H+<����3ƭT�Xn3:��FOC���y�Ó���Ъl6+V��ȥ�X�����@�Q�Zs�qn�~�,��IR�%�J� 璆�T�T sF��/�@6K�E)zB��۪�f5s��E��θ���~�0>J�j���)���U�Fq�+"`|��(�DG�pXwR�/�b�N)~� ��rI�
z��/��C,���^Xi�Lv%}y��~{%�,n��_6*B�m�F�#C|�^���w���Ӯ�:z�u!t�z�_�&��I�W�nQ#�5/s��`�yřv�L��%�N�������{5ɔ���� ���jT[lM!F;�F�h�|o�u�HI��pA{�52�π&���H�wI�n�sbsao�zǮ�/1h���Ý���6C�/�{�k��ݺYqRN4��h}D4��a裴����x��}��т��pG:���m�ê`�%z`�ǅ��)p= ޙ��g���3���Ƹ�#zs�9D�ЮBC�%�y��\%M���*nDsP�E����|!��oV���`��*�b~����;��ǏB��I�ۥ��H�<�x�㔞c�As*��9�������/�ыC3��4�~��QƵХ�!�Pְ3y����R��f5��[��;�qgT/�6����*���Jrֽ}�K��#C�9���6����ֈ�C��/���Ľ;ύXL5oG�`��%�E�k��z� �[9-��|��5`������hP�E��4�����m�a=�Ӈ�_�m�D�b!�'�sx 
�v�D�/�����~־<Z�~9�{K~a)�!��w������ڂԭ���fӭ�Gl֓PY�������20h�5�i��.N|H��x���k=�Y�D��w�x'��𘙏�K�^����iY�? {�,w��b��{�dN��D�@�շ��Y���3%^k���/����f7�?00���q�|��;җ�<z߈�RC���U�=`�����hZ�?�W��d�$�5���������d��z��h��[�,rƋ���P!��<�흃��z)�=���gP�j��F�?��ꥮd턣-�p��/�E�6U����鋅�w?���G�"%�`���>HL�������
1U��@-\VA`�ê��8�%]eV>Nhj��rrӯ��	E��/�c��6ݚh����-ʼ�jJ)�#������9zP-��dR�>�T�| `k�;�b��I�T>�j#_p�)��#�$�w�:ϲ�?{�S=��&J�*O��^y��v��TF��T���TN�8�
c�������Sr�T6u��l�V�KVX7=Z�1��0F�W�J����D��Θ�1���&��$3�7h�N�$7�BjQҒOݱ�ϋ�w��T#�a�.O't@+W��H�	����$�Z+��ƺ���ܵ��,����y�dӸr��CcŪ� h�Α�d�y]g�	L�`%G+��}e�W�^y��4�S�;߽�G�"�6�W;e��cV������>��B�X���M���ԸH�ZJ��� `�XȀ��3���Y�Ya�g%(u�vo����K��5��e�d�3�F�B�<�G8�4����|3�8b�V��sgab�v�e��8T%�|T��-��t��s"EE&EI�����M�B��&�>�*Qt��Y�t#�J������B�Q{?o ���|R�Kp�K'��[H~����&�(�8�Z
Trt.;� ��{�+�]yiϧ�W=�vB1�7�U7ӣ�uTk|E&Q�I���;)�rkn��p�����9/�J�"iX��}�Tz�O�/ڔ�Dxx��ּR����)813E�mj(3�����=k_���~�)�����כ��k�Õ·��������L�a0\)>��BT�s��Tr�?F�H��/,��Ɋ���p��yY:\�L̲]Kk^���G�)Hp>��J5��*H�h�5ok�}A��|�l�S���SA������NH������ :/X��8j�Pc��cVڱ�� �u�u5T3�VQΫ-���H�M�|�=M�-�ߪ+��z�\,���:QJ_�};g��Hz s��z��W"�����!��i*�m�"9d���n�@ǭ����tM+C��|��
r"7�Vf]��<G;��|�wN*�)�����	�`S�p�qs�"\�S��U�]�T$i�s61��P�/��Q��7�n.w�#@} g��٩	���T����T��ո�W�5����z�!1���2�k�x�t!N��BV���aS�ɳ�P����,?3		�4�@�oi>3CY�_���τ��0uK|U/I@e58v���{=P�����������}k(x��kw9��lhX��*W/$�$�v��=.֛8�5���o�ڪEcB"}E�|��=`��5T�}֑�
'�2x��V�ܭ�S��YSuӂi��@k4F���띁���k)�'� �"Ow�ǟ��� N@��E��J���Zz h���D{��<��Jq�BB8tE@�G�i�l��ܐ"��,���֎�_h�GZ/��u���Z1}��$O$�2�Ɣ�N{�Nb���Q�x�b������)Ҽ�x���P���P�}}c�gDM �Z-a�*;�3a�V���!�V�pY��V^S�!@�1R�)��!)�d��{īfҺ��|1jN/���-��X_�o�7�!Ť>�U+�W(o�J�w[5_�'���� �� �t懗� ����*>��$����+V����꺳�B`9+\�0��D6'f��0�X��c6�E`2^c|*�jm��@R֔�:ٯ��=�T��S�e���)�P�"�QH�8��}d��oe���J������$%>X� ƛ`9v�BǞ*���%��ِ���?	)��>��$\��>��&,���x!��s��'쌅�-��/�G<U��~L��K�	$��MМ*I!'��p��hC�t�W	�����M���B���in�Fa9EeN,I9J��6LW:�2j�w�S���mIއ�Cݍ��C��� &@���y#���RV�I��H�q&�Z�_d�Ȗ��>G�6��>eH��)FϫF)���i�@L��.ŕ2��G���n�`��ʮ}c��;�Ħ~�w���L�kqXP��5��K����- �����irZpbm4�	A�\�T��Z�q�[�!}�	Ӓ��3OK�V,��S��s���d4�D�W�[�Ѷ�1��Zn̡rA��	D���KZ����Ŕ�C*u.�ZAQ�b0��mULF�;�9��(JÅjPi"*
=PHӆ��xc��h�����Q�82	�3�x!���y�O(ۯ^´�JQ4��uUr\�T(�KL�{��$(p���=�?z 7T�6����_����#h� ���:p��ȭJԕ[�B�s}*悊gvIYd M�0��Q"�[T<�Na���9J�SEV+v�<��>.�RX�	$9�oe���!�|C�9FY�1e��>\��^�#��%�,Ε��!HRBk������(�˾wO:g�M��~����SH���\-���$�:���<��(�,�Ы7��J:O�+�%���olܰ�P�zN�+�5T:�$y�A��oIe[5��I�B����B^�K*�$6J��_>�Ȕ[n
$��������W)�z�o�ݼZ���w�
����P�<�ₕ	(XA����74
��Q�-���X�i�EE{�uJ��i6�mwyb��J�5R��-)#qu��=�2�W���f���^��B˟��K��.�ܳ���$�][+}���mG�����7m$L��vK�hw�p}o0�k�#X	O{rǪL�ZD(L�*��$hi>R`�}yqmv�["fr�*U��n*�L�Cr�{0-Y��lp�n>��-q:GF�4�j�)�rD�'A��Ay����T�ဴ�i̤�<�d8��>�)��|�S�k��¸S4��)��<BW�M�xY����c�7�\:F�+)!ꨋ���G�H��B�ʝo2�&9cd��J&T@߿*�a�ZJT��ֲ�t]4#�`��{&;+�Ɏ��c�\	�E�t]E����$���2�sR�>�K���a	ؤfL ��L�H>��|S�e���+���PU7���Q�	�R��Z���3Q�q"��jZC�ϧU��)W�=��:��iT�D�J�0�8u �w��z���Pi��-���QH��5�0��Ҙ�G���:"��Սm��M��S�Ӎ	APNbn�MСXl�T��<J1������";�;�
�=�v�	����Y {�ĽX*t����L��k�@�S�<&��P�"�����s�S���͚lr���@y��!�����ډlQ���ή=ʾ}.���]� �q�w�֭���f��R�b��I ��W>��������r��|���!A=\�L%���+ߺt��!����
mV���F�� ��1�1�<��<��|���(��$Km��Ҏ%g1)�t�����6	i�K�I����}�����#����S�<&;%O����n���XV�vL	��R?^��Z�c�R�4|J�O��Z�vT���6�_8�Vy!��;��vrwz}�U�+���/�s���n����2��z0���ґ"t��R�%��ĭ��w}���}jz�@��nz�q�/���2���2��O�8R�Tf�g�X�i�c
�Ӣ�'�kJ"��G��T�o3>�t���k��JWhde��Վ�e���
w�3.ڬ
����b��S�GWki�f$~����u���l�޲6��e�IIT��t�5��uL偤��b�)� ��@�Wt��I�[�4���4���-��y���	RAV	��0Iܷ�/�*�6mUwon�?�O� ���w�"�XjM�Xg��+u-XI��{�08��]��e;���U�����I�9��S�h_����$>ԉVZ�Sn�mN�۩�i��Z�i& L]ɕ����BOYQ�8���X�̵1~���׶��{i鏎׶�����i��9�>Id��\��j�n�%K�x�J���ݞ(��,$�A�d{�� z&~��07D�@K� �0��8�x�}�B�k	)�a��#���u^h��0���kBg�D]�%wg�h��|�N.�x�2�>��T�L�M����ʔ�HI��PRڔ���
RS�(���Z/�����.:���

���ea�C/��l� z7�y�
:y��\uJl�a�ܮ�	�b^��	�.Y�ɑ�=�Ap�g��� �?]x�����nsED����/�� ��pڴ�*�S�T�Tp�*�1�_<\�9�r�s�M���nǀ3�  $ٞ�@uHV�r�ti�����P�M4Vd��N�9S������B�ił�����T��4[�	��t4��b�8�*bgr��yG���?I�hG Ɇz�K)&�-� d�̄j+���"n��AR���d % IdMV��R��m$�S�ӑ�^��˖a�[�N�����lZ�@Q��;�����U�'�CaG�,�!:p߸}	�)�$q�8��@p�7&���!H�.G������e*l�F,�z7�� ����8d�I��]=�lq��`�-2����b�д6�jl�\��`N�9a�H$y�󬙶d��� ��mhD���+���A�I
�g�P��O<�V��"I��*wх�s��rU����F4!��r�Vv�SBq���k���W/E�TO$"��'
u����2�9�m�H�ms)�#�5��b��]0^yx�s���8��9����V�f��8�wX�y�q�5-U�H&Z��7��e�\�YJ�\��1oôAn/�K�n�.f�v����Ӄ	M��R��Y��-��ڊ�&F [M�G�f	���*�c�4ߦ=n��k���b۱.�N[��wJ?D[��
z 6t�����9+N��y!��aD���8��>B<gwT8�J}�ʻ�lU6�C[wH�P�ث(N'SB�;m���)����kf�-6�c��ZP�EmJv!@��z��7M�#L��-�q�,�W��Zgk��4B����p��<�������7���G1eC�ڢڗ}�	��uT1K�/�3�	��WP�/J�������,v��#��z,��Oz!���	�#ūd�Ix*Z���������e)��������>#��鍝��ԹhŽ�F/�(�͹�`���7V�*Y�U$��f�>w��^h|F];�xlhH��j���L̂՝W #����#�#�v=��ac�6�
�DZ����9?UP��Rv�Z� t*�G�h ~�DǏ��1� �T�'����i���-)]C �e��"�(�!Մ���&\� ���o\��*h�+O�&X}y����u�yБy��=�$�3�
}5g���E�2�x/7T�%��0�Ȟ!��ʵ���u�#
��ڏ��|D}W>����y����k�_凕ght��ѳ����#�qwz����ލ�$)�a+Б�
�b�bް脊��sgԵ3r�L�dH]��E�Նd=�C����~����\M%��/>��{��*P��u�x�|�� rJ;�Lcؠ���d>�?J��K�B�P�$5���q)*i2��»Ƃ4���9k{�Kn�p���&`��gU`� 8�r,�i߁�#�� ^b��0�!>��.LWwZ�Fխ�9���O �k��Ϫ����04��q�g���^�{�)Jwî����J�
���k��F���d�mI���@N�k;�d�h@B-�ꂣ<��x��%�<٣b��/�|�{@���g,JQ�E�����f�U��xvlCy�_���VZ��I��l����ا��
� !n&m�-�nĎGv�J�M;����+%RHai�:�\�"��6���IH�[�-�J��%-�串�������P�GZ�ͣ�D�V�4̦�$�|-I�-R����o,atM9�����:M�Fɳ���>軚���@���ՠgI��dMC2�&r�h��p��qz�q�1L�j����gu𷜵n(�\'p׭-�t�W��!RG�'D��	��o�~葿��j��dN���C]�E�KO��^��g�Ӳ�nʗGYj�'���ݠ�+���T>��JUU����pK�[2�#�*iU�+�O�^в��Z��<wUB��B^�X�q��
��ӝo������ЗV�EK2� ��1�q$�MV�Fņ�[�LVV(�0qS�pU��<��ūV���#-���IG
�&��qb�'w%��}��a�f _-�f0V�C�x[Bj�LS/��ƭ���0��*A��������S!��<��ړÊY;Ǽ�6�e��� (��3c�� oLw����t�;b�e��_���&L��Q6y :�J�����TYuGZ�䙅C� ����3�� fD2É���������4��a&��5O��#��z���ٹ`S=��iI�����8.vh-*��ޏ��:�����#�����W�b��/�Z$w��I �;���]M�����	[ڈB�ʸ@�KC�b5\A�P�b��{�[~W=L��*��<4��t�%I�V�a��8�Bׇ�y[�bտ���('�)��U� 樔��.�V�u��-�9�QK�l���z�ꨨ��B���}v"�З���4�k��?��|�se�o��lH@'��U�!ǖJ���ћ+~���r��#+uA	��%�ĵ�4eqN�w�p*-���� 1�w�?���%��~*�mX��TRsJ0��S��DZbj3:a���8�"�L�֊�&�NN�a	�.7POٸ�D��Úʱ
�14-�p���4o����%T� L�3��V��$���-�Yn��2�r�O���m�-GU����<�WWh!�Bhi)q[�S,8�r��8	��	�dz.u��*n�'��q�2jU#
���yc0���p���uրy�FXc
�⤰o	�HƔ����jL�X�Y�(�i��J��x��pEE:'��
S;�"�*���h#��<�b�Q~LѵZ
�S)&��Z���Ӌ��
R�J�d;�1��v�*X2	!!#�&��T�N��׻�
�p�Hsfx/�	'囵GB|`cU(�j�Cu�6�ȶ���;D����Y��
��9$B^�*��n��	<��i�p�$�<�� 39���8mB���{��eUV�)�$5��)'
��_���,A �%�d��'��ʖt���#��\u�2u�� ���H�8��2f�zx5b�� c�ei
m�=��d�����iA�*Y�0��S7�/`��M���;��*d_`�'�92���;t�Z��[�ou��� X���?�<�D,$�e���b�1�:cQjG���.!g�N��CI�~����T�X��Ɏ�����f_mM�Z�BS��=:�D�"��cw�1Gd/�p�-)&|]�<�p/�l���I�uO,R��{���},1T����bI��$9�r<-�g��)n�/)�(�X�h2��	M�z�#������nhw�Ϲ)%� l]ŗ��N��	��ų'�-y�0��l1O���X���P�h+c������l=Xڋv�gy��%=yO��"���	�_x��!;[n�2�c��ۊ)XH�2�e�+��(� ��D4����HI�R�FC#m����!(L)+I�����O�����Q'�X͉󘲖��4�s��ԃ���ç��bIا}-��I��Ѓ����% �4��ɴP��l�މm6*��Y�u=I��l����?��x�$�$�o��$�ݒg�a��<%/-���y�Z�A̫8Fr��O�=a����v�� �<�.^��d��� ��DȚTG�1֊d��^C��_>[����9����kp�[W끥1��s[`�I�H�̨��!�=4���*
Hi:sŻ�>�%r$Ì�@ⵕ�٧	��'1�0�����J��GW�j���h\�l�Ɖ�\
������o.�l�� �e7�Z7ߨ�/G�21��,>��l��������W�V5�dV	� 9Yd���A<������#���5tGf{�j��������
�+���Y.܅ ��Z,0�'ℒ��.��K̬���T#�+�=���tBMK�wWi�͊�n�)6Glw�
M[�6wߨ�+|��ԭ%iD�|J�D�*8�%�����?�}1�P(?��L�akm�.M-�4K��
OL���H.�rr۴�>�=n��쫦,{'������7�}0i�@�8���JZa�]�\� �Yh�M����t�J~Q���ֿՂ�O�Z ���+X���� TRҫf�>�
�L���H��� � �:��|�ŨY��q]0���V����̛B��)q�`F�x �I'���m%j��1����
ާq���K������yFJ��L8�F'C��Z�cq̜Fv���ƏXC�bT�KL�j0�V$�I�?�-�@BXA��9ϊ��J>���m�!ǋ�e-�q�8�B�>�˚V��M�X$'��w�W�Bp��F���*C���&6t���y�wɉ�Y�Q���>��o
��,a�C���H꫐�Q\�>��~ʣ�9�>�£�;�*;;�º"_.�j+�>�¢����i)#�ʖa3�22��H�#}�"sø�b_Dz0��8ZKxV@�b�>�:�8�&z	�N�&'�7�6�#����g�w��4��E�K0̐t��]�u?��m&�f��&s�nr�+9���1xW�TI:��z�f�Hq���ck�1�[����UGgk�}1�Z�}1�Y�}1��]1�g�_�Vy�V}����OLH�~�����iI�D��7O���� �F钬*rz�xN"s�f�Ȗ�;T���`�Z�b�0���TuZAW���f_n&�(���0R��`�d�E�pG��� �氃�\@j�I\ЫK	��$h߅��6�#�a80��MC��TǬs�xJ�O����Ց�]�~e(L{�8�ޔ{���>�@���%ͩ0TR$H��wp�����"�Rm���T��ga���� c����T��@�"֯X�QOJ�f�z����½�ŧՄ�C
��>-W���*��yi�Z���G\r�p'
Ұo�+T�fd���q2�bb/YwTčRA�f<���qZ�ď[Lu����3��s����͘N9[�
G�2�ƒz�1��{�l_.H\�q�z#�<T7�u�H���Yi�1�G�|dr��)��E���G_�E��ӼDb�OZ��Q�l���I�p�y|\���Jc��&f�-*�9�j
�#C�﴾�a���U�Ԑ���	�Y����w��İJ,�%l+��N�h� �J'�{���q<R$��Q"����b{E[|���F ��j�c�s�m��*3�=(�t��Luc��lu#��X���0�b��!���yFD���M�ڕ���~N��k�t@Bu�p��%L& D�]<6E���2���,�7�<�����6nS{*�d�FC��Yp��d���CBE���9��#~s��U��7Tv[��cV-i&���H����CJ�Yg�'� RR�X��'vϫ���I��Ze��ˆȱ^X�������T�:|Z�.q�C���gN�aq��59���EB�5R���T�-�(GϿ�B��ف�~IN/��X\��W�آ#�>c]����)�d���%	�J'�Ĝ���QiV�ՋF\A���&��3Y�<	U;�k��e8��\P�L�՘��r��_��PRXI���'�g��Z8�C>X�=S�i���f=A���U8���3w�-�9��-#��d���?�z��`����2�y�����"�� ����0��������������Tx)�t���Gh\�E����p���c�9[i&,i1ci�T��pA�j��|�+�3Q�N�֓�
N�)��Ǩ?ds��Uw[`!#��H���w���c!8��4��,w��&������Ј]Wv���Y���^�T~���D��O�-9��-�6�yT�R�$��;�b�@5� ��ŰXT(�����Q�!�_HR�ʅ2I������RZ��sV��E��S��e�#/Ϫ9�ds��SH�Tu���q<�f��@߻qRs�W�`3L�nJz$4�nw�f7ҠR�D�V�M���.(��vx6�Q����1�ё��5�pq�8f#���_����8<[�oY�F��YR��<F�w�~���!�S�+��ڊ.RL� w�� zj]����SceD�hL��B�G7���s�*�H�[A�膈N�������T�ƪ��_DZ$s�W9��!�n��>�R��肥(�f�(�n�Ԩ뭩7�3�ȴ��qe�68H��6�+�U�Si��E����ʮ_qx�ӰgRG���jQR���.��|��}Ӓm	��yb��`N*] �W=�E�vK��m-`^R	揀簨���a]�Ɩ�tԒ9��z�'�xv�	�y��9c�\��8��x�m��Y9₥��I�)�d�VH�G@�m�ǻJJqX�����)�?e�����<�J~��%8ox�'K��E�t]������R+^�8؞�G��X������cB���DLeOwP,�SS�$��fJ�x���N3 ���H��hk�54R嶦�4nZ�G7��)�E�E��m�v^���Q�#
N)�(V����䧭#.KRJ���N�]}X��@��I�Ɋ����14�x�4A��8��Ú�^R25,���Ŗ��.
O��2)P&PUu��xcj����]8'�L>���*1MkZ2HC�ۅ��!��
R��<���em�P�	kz0I�0��C|��b��1~H��O����[��Q�珆��H�#�!��(W��l�l^�8̡�e����b�lW������bI*F٩2Ju�R�u��G� ȲyFJ|ھs@b O�mB���sT��%]2�4����]	M"��a�����	�v��k��qr��"��oꌮٙ��!�g�Cg�� h�.6Is�%f�/���4@YIT�v��Q(N���M��6�$��N������˅*It �ᆝt� �f�:�a	[���L�+nÃ~���:1g�YZ�ժA�a�U�{%<����j�6�j��U�uv�$%�L�H (M:�_n����T'A7�u�cmDIzd�'����4��D�_X	O�=ڥ��f"��P6�4��XM��V�%��E 
8��b���o���q!�!6qdo�'��[|�]f�T��^H�_�G��I��G
��#����� U�k������S�����M�T�i���[UL?ԋk)���ܦ;m?������������"�#����j���}$f�C�� ���pbmN�(i�Х�,���E�h��9��A��#�&l��� ݋OF8<��d4.ZL'��S�.~]Ө:�@�@�\lf�
���p9���w�s�^r�	�%�n�d�!��BW�`P @Yl6ۍ�NJn�'iᇆ��n�8�;�m��xpܫ�X��=T�?�J�R~�9��[�p�A�;�d�{����˄�o쒟,$g-��D--�S�FxJ��}8>�8�'g���$2�LWi��J0�U�p���*�/�:�(qp�xzgD�J�T�(NXb�Ր�AN�P�=0�ڥJ�"d�|�U���j�����}�A�)�����T0Л�)�S4��*�p�E`WSl�	�'<H�����#�I�ғ�����hl��1H�	��7��w��Vڀ�
WL���xj���&�~���������l*ZN�z�z���C�����6�*�R8S� � �5�S���`�B�6���V)�i�.�ZF�!ɄOZW�u���)�^�nL.RT�ֺ�r�(� n��&W_-0���1'�e)�P�H3%G|�(si�|'�ڭi�r�D>��l�L�5�Jt9� �L�8�ߖ/k:��TB�Ư}��L��'Ih��иj�*��q�'
R�Ӑ���ж'����T���P�K%R��\O�¢�1*i6$�1�!�����D{M�a�eE�,C>|��w�iV��IN2p�;� ��c�=��}0�wU)�u�WYĬ:Y�>	<#�P���{`�l��.���y��ioӵrNi��;�����\�;NmL�e��<���t�9��f��i�
�ԧ*\�Q���:��f��BU�g�7➮��/����2ft�q��4��Z"���������:�T�*V�����)����-袩�X] �i�J���P��ӭ�5�Ft����Y��^��sfWؗUA���y�u�J��_4%ƔP�mJ�|���e�"ßxy����U1�:0�YR�)*���_v��^�6�n�o�jN�
K�\_X�(ާ
����T3��p�m.-�	��'��aUNS>��j�'S,1��
4�JVi[Ӓ���M��H�y��XTj��|��-]��	i,�5N�"���P�ӧ%B�j��T�&d�ӧ�(=Ut�;��zE	 p��Ʌ������V8ٚf';�.6�s����7L����6x/F.p�F'd�G���bC$�E���E�|:�F���1��g�1cK ��`��=��&>�ɏ���m�Q2%�z'�^()P�o�;I����jW�"ڕ�";J�v������R�ڕ	LF���X'�(�$L�y6����� �3ڋ����1������� �]1ٓ�ʈ��Gekَ�ײ#�5���{">>Ȏ�߲#�7��M��#���h�Du��G ��䋢�(�,�p�  1x�|[���ķS�n%� �������/� �o�� ?!� H�K�������� R� �����NgF΃)�9�M��S`�߼����y?n'�?�Q��i���>��J.wT�0��>@*ʜR�Ԭ���J���*��	WYhnX�5G�IT����>M㥀��� \�b���H9&H�0y� {���P/e+1	a���)�a
��ry�A<��� �S����]x����O��{�k���1M	;�)������g�*�����_����R��«|����O�����<L��f	i��}��($�&o�ܷF@��*?��+Қ-@On�M�U+�����P�Wn Չ0][�� ���
n�5�-D����.W|����`-״�V�r�?Hl�"����Z�ߢ�5��a7E�KfY~H����S�>�r�n����J�l�S�Вr�"/(�ocr��+��(�v��94@4�EߒB��!�8\�QƧ*-����$#I��� Q��� ��4	q$�X����wAS�:{Qx;�1B\�� R�5uȎ��`T��F��v��	��G0�~ӨؾQ�콌�+��BĶǴ.����d;���5�epU����y��� -{;�Ж쏥��FTx������ߦ�.�fuB��ݪB� O��e���I����s>)U���U�G�h�Xt�u��Ս���3-�x���C)�BO���Q)��pb1_R�v6Tg��<�ۂe�\Ga��h3_������?f~&d�:j�����X�Ip9� ���-�ʍj�?�6�[���Q��������I�Y��M>�i}8�����SuY�]���;�b���+�S����p���~H pD�j`.}�O�l�Ƴ1����ve�\C_f2�"pCu�H��|��f��r��y�� �\�L��	 kWk���FNy��V��`������UF�n5�)M�Yd̫�������F�����f��F�8F�J��z���/5���M�Q�	T�7��{*���e��f����T�^�����'�ԇ��x1l�L� C�_A/(X���ڥ2��w�Nؕ��>��rf��u�<9�UƢ�TA���T�E~U>B��cL�U�,�(�]Ԫ���2U�%�L~&2�S:%�9��u���1�I�g٘�̨=�d;�����-	�),�Y+����Uu��y"F�����{��:#���@�vŞ��q_�++żMy-r���LjU`�Yo�X�$9A����L�� �-c�������:L�}w��������$?`�9��|�Y��pT��H(x-fD���O��﷩�au^�,��iB
��i{�7����~�"��Gw~�� �iM����[C<�f�|rW|�29ʏu��dzK(�����4�;��X�Z*Y���^�Y�s�H�>a�����ٽC���������=����BXR�]�5������{�*��ӷ9�"	�w#�"`�5��ݰdf�?��6,~bo�m���㋁C���bPg]���>iswy�"�";�T0ױ>�.�̼ |�c�v9����|�^7Ya��vw�� h�#�'N�������y�١����,�ʽvDC�R�g�YF_ C,�TZ4>�������"��ffa'��ľ��J ����C�8�Y� �S['���?���;	4,�g�b,Ug(=�2G'��������F �2)�} �{��:�Xc��G�>�%F��	�����\噀q�ʊ��r&��1b��t���
��t\���*��\���'L��jŧĨ|��<ec(s�2�ý��߃��cvUJ���9�����{	|��h1����KQ���W�[B(�v �����Lj�j�����ߤ��=�:2Ǒ��],�^Y��d�J�j��2�}���U�|"��x�(JKkS���N��qg��F�R�J��d�np5VD�#
ޟ9�&�|��F�GUY�q��]��"�C�����s;�ii.�q��w%��gw��AB|σ��(0���q�,o�+�1���<�E�$� hOn�w�����M~Tf{��ac�=�_�!1�)�
���0�
�K�o˟m̝��\FNH��A��Ϣ������qqg�l�9!�j�WY%��Ͼ���(	[&�bAg��{���./BƎ���?���(�fhS%������r��w,�>'{��_�jy�\�4��\Ŭ,~�>�7S�,ᯩ�rZa��Y�~���b�-Ф�lH�����;(�8�p"�W؉7UO�50��@�d���l@��T�;�>�J]ݑ��qD`�JǱ�Ur��S��iu�A����DR�+�@ �\�j9uٙ�6|�y@�V'�s~ �.i�,�i�x��L�ܹocq��著���g�^sP8#�y�^�楱���_C� _	����@��6;C�q��_jf{�>���O�*��H�0"ea�	��1"pN��%�c�b�.�%W�+7ét����X��o��UjQ8Nnk �碥Je\�iO�8T�UJ�60�����^��`��?
΅|���8�(�UHR=�r��l���P����Wy�0ҴB��8�)j����tO�d[3��v�Ux������)���x� mN�R��ǿJ���:�ݵ�y�#`rf~���uqGީB�q���N�S�	ġ�S��Po�N�|ըb�s��5B�׌�a�p�Ehn�'�����\�ܴ�8��Y��(�*f��t%�\q���,7�O��R�3}b[\�h]�?�|10��I�RhB��:��}7
�E|W�TYk��(���rNܗ�. E�Ýo��uпF=����3ۣb<��RR������JK�.\Y��������Us�l�9��6�W;"�h?��%xAh�J�y�R�q�BT�S���e���i4��%,M��l��s�O,V\Y);��)z�4�*�ޖ�����=%�I�I�I�s�Qe�x}��[�ӟ����0YEJ�	Sc≑�8Ǐ;RD'����s]�ٺ�t�y|�D2c������z7QL��\:�鉆�������-�qj�&�2�瞠r̮�Eؙ�����[�*W�5}����5��|5�iC��D���p�|x�TҚ���͜����V�|�W�F��}���x$ ��YGyR�Lt0�F�Eô�P�������$��eY<)���H�}�VVi�W���iA��(�rs/�[��+䃆��������,��ۥB���n��w��(�!=�Zp~C�~��6��Y�{0��h�J�*vՋf\8]� E�J�auaķvߙJDj&�e�v��R�J%@d��фM%+'��fecpݩ��au��V\6���X��5j�baų���'���?�
� �� b�Y�u���*K� ��C��B����0Q�� �0\~�2i��*� �l-v��&��E�+(�4��!h��.�i������ް8��cB�No��zS*; ������_�~:���B���y�eJ�]y;O�{��Y_tL����ui܄(�"a�0�׀�g�y�92�TC6۴x>�SG�C�� ��S�� S��̿t�
	�ǔ=�]�f ����K���៰�M�J���Ws:��d����O,ǒ`�6�_۴�����ycJ��O��8�uy���y�����lH�0W2�]	"&i���.X�";�`�$�_R8�(J�����p���G�\;y����S���J�v�������+}VhYD�b��/<�3�NV�������,��h��טf��B�$� �kd~�b��Y5�4X^�j��9��9(S�왵��`@�%�x_����^N7��*� ���_`�q���A�\`�l[!�1����^]/�����"m)+�8��߉������o�{�Hd�̡x�Hv���ID��ۣ��3�Y�EJ�����9O�!Ӭ)�J�K��y�+�R}g]�UX��pf��EB����[�
���T*M���7J��?��A�?��� C�?�^���>K?y2��{t�?v3e�8N��> 9g��k+���Wa�w�J^�L0�+q4&B8�\;2��zF���i���\|�Y�Jy��>x$n�MKEÇ�p����׽��!��L[�eմ6��ʸ�/c܁����<|�=�so�eV��`{��Y����,����L&�Q�@i�@<�W*�!��d�����U�]d�`+��Y�8�E�W��4��3K5���,_�{/��$մh}��y2��ɞL
@�[h*c6')P-/'vk�� 5�.G�@���Ol�1!m'�B�f��C���Fj6\���==��n��iR׼y4yw���X�tHs�%c* �4T�'3���crm�p�ok�R1��K���L
�9bN���,����z�(Qx\f�[oo�	�x?CG������rm~���2�b(�iK��Eo��JDQur��2YZ��9��	�9Y��.5n�fQ=��F^��-��eӧ\��璌2GD
�����i6��x�A:��R�7��iB�~�5D&~��?}����K�����=�L�����Kx�%��pU�"=����aWy�-hTpF���	��@?��»n��sխW/����*u�.�ÉB@�b���EjF��nר�џ֜|�Y?�U�$r�A�6��G�q���_A�,O���r㾏�>�P�u�Svr�!��n��ly!���o�M}e2��h�ÈNZ9�&U�iP���R�u�/9:P�xQ��~4�缫�^��;�FJ��{N�m��ǩ0��#ݩ�(G��a?�Fg-��CP�ᣴ��(s����~p��M�(6�����Hi(���Bh���2�<"Ph m�!>��g�� $�ўvT^G?�A��(`\��⢨g�kܳ�?�.`�/mJ��T��-�d��[Gq���u@R����.�4�)x�*�md-�q}�2�� ^*}�mW�;�%�U�؏�k[�S5�[���M�IO����jڡ� ����7�+4�_T�^w3cxʌZ��X�]	�g�>d_����e���]��H
��ɛ��d�׎H����eP]Q��ypww�w8@pwww��܂��[pwwwwg��'�[Sj}��W�V�����U�����38E;�� �~��P
^�YEx倃�!Zrt6�L����8Ʉ�Mj�b(�q�8a1�����tdŻ�r*��$��!���|��1��}��(��2��h�G���n�k�.ݐ����c�Z�{�a�[y!	=��8���s�ڪ��L?9�d.&;$Y�%z�>v �y�O.o1�}G;s
!l��d����_gn�6;Uy�y!R�.��18�f(�ؙ��m��*e#�K�8�)���"�s�*b
�`8'or��}E��[S��V��� 5t��LО�3��s�քpT,�GF4Q���<f �\.8P���h�)q��y��y���t�q���_��tD���v������2�%Fm!�3eX�3 �V�0��z���hgyb�J��Nt��xm���v��Bi�<;�S-2�ם��;Q�BO1�o��u��T��"tM�c���+����՞D��f����h�+��������c���V�n���mپ��[�9ɴ�P`��W��̈"J�a8�	TG�:�s���JxdCe�u�k�ն�8����&�`p�v�BרH:m��[uQ��OB�3J�t�&Z]���;n\m��	�xk|�l?a%�-�(�����!ZS�����ZJ|�AI+�B��{)��z� ���z��h}��0s�j�����K6-��9�ĒJ�^�4H�jv�჋�<��2j�臶,܌�S1�,�{��U�{�������.w��=�
X��8,5@VPG}17a�����	v�o`�:�/c����[�7usQ�wM�cC��$�
��)��<��v��#�g�A���&�V�
��M�7�%~�+gk�g�������e���VM;�G |Y�X|�ڭt筄��݊��pt��k�L�= ��̐�6���ʹ�P,��s,������$���խ�J�>����N�=C�&�A�ϧ�ub�>l�2?�����\YtUK��~d�@X��*�7��׸ֽ���?�؅-!ֻ��`� �u�|9��QS�t�k| ���v����I9dU��H�r�]�^��Nr��rQ��x�7 '�"���m]�1�;��{a���V�r��L��ۥ�.E@��K��-;l$��:h�t�r�Р�#��S�^��T�j�\$�i8�l��ś�
��F����
���g�jx|?���{2Q��_�6vB �u�Dn�������N H�h�M���Ydߖ���,����c�.��z�D�ev���p�Ӎ������ـ1��N����I�xW�L�s��K��cT�E�E��.�PZ�U�
�����d�a�쌡�,��d��@�Y�_�]���ī���a��`-��
y��%xM<c��*;�%�r_�Xҵ҂��`������{,Aἷ�飹GO>��u���V�'�M�?��Iu+���D�E|#z�9`�K���%��I�Ҹ�F�l#<�r�ia,����q}��E�%���%��j�A���$��`��,`=�˷��W�%p[���C�S���j��	�Uw!v��tJ�8j<%�<�z���r���P�blR�L|1'f�M/�:�%�5$X����O��� v{^�A��r�����h�<�5vN���1��e$�� ̢���U�q+�ѕ��7���;
f!�k�� �*Ÿ��cz`�SÕ����K���g������r�%N27����/��|S�m����x��s�CE��t#�ߵ¯�T��B�R�JE��2B�{]�P���\ʛ`��+�����p�1��x��x"u5?	U*p(�V�w$�<�^2u�oJ˯�i��RV0�����㫋��O�]I���4�Q�R��p�o�CB2�����qW��s�㧛�7$g;���9ؒ�S�@Ԛ�j-7�1Z�����A���n/�
��=�amz}���xb��s$��2���UHd�9����^�F|Ao���Bi0[��"�H�x��"�qi�j�!o7��X�`c��q�A^�����%��sn�-�p�s4k$����a���P��q�qd��S� �Bq^[����yN�B�b�eW���B��B=�o4������Y�]Ho�>CR��B��奠���Y�A���u�|E�(�
�ק�Y�o�|�<Q�p�L��*$B��(F��o��v����HV��dV?{����P��Ar�9��Ϣ�cK�#P]�O��a�zu��yxz����a�ߐ�t��@V�}���<��i:�E
���|��O�x;28�.C@����zÀ`�T?v�=�,��b	T�Z��OjA�L�����C}��Hz鯒pd:�!�U��tè5{Lq���B"�fW\�_=ϑ]��Z��T�{��]����Z�ǩFU�A�+&�P�WU,�S�����J��҆�G������~�g�d�@?����1��V,
��"�k�� �jY�޾&E>_���t"%�����X���i{쏋��{�)sx{����R�� Jg Z3W���D���I9n%H��M��!��u��JKw*�!M�������ёK��1���K(jl����c�~5%]`��2yL�+��?���������йIsƾGf��~ƾ�A���`.\u&J�W �~]j������D�[/|�q�mH����u?����VG�1^�iH��N5��>�D�"w?=d��H{UM������*_�I,1/��΃G���y��u���l~�#�^~iN%��:��.c�ו×_����jE�w3R�� di�^i&UbD'������ag��$B�#�n��d��!��o�J���r�;b�tg�gDU�i1QBJKC�wp�E���照�YO��'G�x���� �V�1o.D_���~���k\�i�~���:= 
ZEP�"4��*��|�,ށG�W�ڋ#2y�n#
=����ؤ��n���/^Q۹�p���w*�Hx8��^u�Վ�&�Zӛ�������!d�8���oĶi�+���Z���C���]~�	��V�M!Ko��>ȳ���ϫrܿ�>���
�� �`C����V�MBN�br�x�۩��dP��M0]o�c�;���9��p��Z+`v}��k�
p!����7�D���W�ؚ4;�\���΂"�;��;[ut�q�i���Vv���[��R\�B���g���A��͆�ƂQj���JH���˚�Q�{Nj!�v$j:]gڣ2U�m���f[�r�1��34�fm�����i'o���-9�1��ʋ��O�%,O�� Y]tpYju�5"`Ni\i�h���2����m�ⴍ\��s@��4�Ef��f�_�n���(y ��#���wRP3+��	P�,�/���9_�
�g"����z���hH���3���^��+Yx����U�8�γ�I����3(�w�G>�{�sYjv���0�3���˃%�pF=�L�n,9��+���$�6�zj��:��e��.a")�I��7b�TxZw*+qt�ftO?����K�ܫ�M�,�P���;�80�kŁ�G����b�]1T�ͻ�,��uZ[��A�>͓sO��DYZ�[=�0.�^7�9��H�~ �1j�A����})'���mE;f%R_����O��5�l{o��wК�t��p�	�n����ֱ\��z�;��C���mi�ݰgx�ݏ
v��A����\��RP��q�w7Ȭ��˚4���vl2�M�o�oI�#���@����]��S	� ���!�M~��z|'�ꋛ�\C�ŒP� F]?[�+�4,��-;���0����RH:2��!߱W�pF�ܞ��h�����|�Ԋv�/
P���szlּz�~E�C��7��\�L�T�II��SFBo�T�a�
��pIR�����W����)�=0���OIa���4�qPE�L��H����Q�s�2�1��j0jµ�q��I����e����d���9���y��C��'�`o�(.p�q���|,����ʺ���Ls��-��X虹^�kr���4��5�X}%�D��H�zP�s�"jhY��H�`|Z�`ѣ�+�L�' �:@��@��m2	�M� [�V����œ*�`Å[�E���|�t���$�k��W� ���Z����f�^�A�dĮ��K�� �0��n�&���-�@U�Ł9v�߇�?���K13FG�,�[��45�:��k�v�����W��b����D
�5�ӎu��sE��Mqn{��+�2�}$���C�P��B&*�Ậd��o�>�o3���.a��@�E�ʴˍ�p�g��a�}�E���E��J�Z~a4��&��`Z��,,;�f��Vac�S�`�N��X增Ѣ��0�_���ƣ��O�,���+�(O�_H�T"N����}
_tP��K~+{�ΐ>L)Ec�M����{!�UP�}�sR+(�p��p����)�ټj���h"�OTb��MZi�"��h���P��j�v���21��C����;���>.OwA�����ǟ�5s���L5�֧W�c�K��7)�ԣeP_7����z}@SWf��b��HH�)�R/��8�4��3d�+�%����/e���׳;ǻĭ7�կZ����3��s��7�}�+�p+���f�w�*oxQ�����~��,����q-ożW�ޤ{?> � �
���C>)��^3�o���
G�郓�E�EUF1riǱ�p{t�x�Mv���M�4�(�� �\u�b��ha�8�5��:�'&��v��s#*)��\��
c�,_�|�h�4�+_掴�U#ٰ�ٞU���o&zR�iD�stJ]��?�D���`���P��wK�Ϯ}I��]���	"w�iǱ-˓ّ~)��c?9��#L�ct�]�*��u{�)�{Ck>$�s%�)�w%����=r-$�ށ�`�Ԧ�٭;P���ib_����
iN��>>�g&��F�$���4�pЅ%8[ȿ5�#ê&�a�?u�&�A-�-�Ĉ�;B��޸��Yd��Ov����0���oj5�لL9�b����.�eW9��ܛ�7����>
��Fx���3ÊYk�s��L�5�u��p��@�f�a�X͋�$�I xe;����)����
��􄆒h淽�&�s[���K����j�u�{�LDu�3�/:��;{['����jBTYBې�V��}*0"ϴi�	�r%\Ԗ�@.oJ��j�Ū�c4�V�V}����ŮiP��XcO�r�1��-Nb�2K$�*iSd��Ur�!\�r2�Q+.��=�	�+��\5��Ǣ�$��`�q2d.j>�]M~��!Ͳ�8�S~�0��ٺ�Ć��u����e�P�GBz�u�����67�e�fO@��f3����g�b�0�"~�Ld������n̕�����򜛁�6��X�ح�R�Z�k�w	���9��Lז5n?�H��!�(��̛\�P���vE,�b���7�~r�U\w���J��b�S�dz!��Siq�GX�B��H;H�>���������^���$�8�5�x�y2P��A������O|HA��uT|^ �����..D�~��yl̰�<u��'�h��z��F"��1R����'��OL��n��bGc�j_4.|�8����q�h�|�(��1�Q���rz���j���s�ׄ
G;jz�����岠��tB�o+e:�:��<���A���>���.���B���ͣ��m��05od'��gѪ�9h�i�����yK"ȐjB�φo�vL�w��T������n�(k�}H���Qb�+�'����<9v���uإ�A��a�%�7���!����o�i��XVʹ�ܮ`5���Y��t�,ݯQ��`���F�m���s^Ѿ�4F+�6�=�� 1�$X����Ul�OȺ�҈�W?g�
����bw%���{����u�(�Nr��|Ǥ�0Y1>g7�;,ߦ�?�"tA�x}�@F��Y�_a��+����}l���j������v�H6M'=��0b3O[Hf)&�/g>�;�M_���ŉ%��t��^��D�mB���y[��)�S�d�����͑����_�8i!-B���Y��S|M�ݻ���K�>߰����K������s���;I�h�Ջs*�
�1_�g{E�������"��w�c�5���������ܶ5���U<ܸ��ԀNQ���תY`�67WD�zn���E*�e����w��н�Rk�u���lg���f��=)&�]<���y������ꉝta˭B5Ot�-��SC�A������\8��~i�B[d>�U��p˗<�Bc��]p��	k��}OR�J�v_�R�����%����{V��6��(u\-��]%��s<m�Uc����q>tV{�I�p\�dЅ=�"�.}e�����՟�6pv@�?�}��ϓ�������p�>�a/~��v�=�"�cH}[�M��K���r"��� j�����P�]�m�/,g����p��;�M�*EJTB L���MD�8��勔��]��bm�,h0GrW�n�m���G�b%��#� ���h8<O��>W$h�z�L5�6�3a)@���ݵz� U�w$��ll
�xH��d�H�Aݾ�oԮ�
������>�A�8�p��n�_$���w=��{���gʬ�|K���p���3�>?:�[/fq�? ��1b�t�#\1��=_�+�D�TV����<x�<�.kh����y7
i5#�V<����lQ9���A9�$�ӒI$r��$�<V��� 	gSJ��)�©�=�?���ҭӨ��\s�S+���У���=�p$`lZ�E%ޖ����2v���cxf�`�>���SrZ�^��c����
ئ�'+����y0#��q�b�{���PU5@^���0�핼��x���j�'4��'J�އ�F�?MG��A���q!W<�Uf�=�h���~p�M	�M�V59��P��������2��,�/�	{/�	ٞA*�✀U�,d�Su�zo'up���Ф)��U�9y�5�%#%�S;\�uҤ�4�o��8�t�S���3[3��F�sȭ*�{iE@Rd\/Nb�N �p�D���p����X@�F]'O�x���˳���yݸ���~84���(Oc`}@Z��Ʀ��j�پ�F�b�Aߑ��.g�k}�)�1�t����������7̚T�)���s��]���G�G��Я����B|=� �s��W�M`�S/����E]?ŷծlAHi��cG�<���}{~o����M)/�G`�5wb;�5��J��������s� ��2"�ҵ��7yn~ 6|ꐈ�^|%> 8���N��6T\�8@�8��n, �,=�����
�A5} �D;s۽X+������,���zp�xjQ�G��罚|E�^eF_�30QӦ���֚�4���ާ��p�L�8U{�,�En=	e.��5f�8�Q�xt�W�R�E-��8���57&�h_��!�P���)��Ce��Y5����6a�x�Elo�36��\��y1]�ad[���KRղ�E����U 2J+5��>��ټt���w#�s����5������|���J��
$F�Se��Q��nv��7��*ٲ�<,\a�Vw֊|���H��?�hS���L��ZO��N+�5����6��������KX�+�wHq�j�舏��3-�4�"�gg������|G[�SkGڦΘ 6IZ�Mr�(f2`��@�%�8��b�$�0#<s��z���w,�'4��c�p�O�������BE�k���̙�C��j�ɇ�46F��~$`��Ν�?k�0��sN{*�$
�����D���O�Rc�ɞ��/� ~ �t>sB 5B���
���0�������Sa½� ��Ɂ�%��> �{#IW�洺w�^d���>���9�|��@b'�@Q4�1M=�ٲC�cZ�o�E	��ߙ�U�'���y��Ŷ�2Ų���n�G��Ħ�k/�m��E	��"�E����q�a,f��y��y������l�H!�����K�2��t6n�8p�]�a���9����%K�.>P��J��4�Z�<2�=ԏ| �T�	4�>�$z�@��%��9�@��6驊|�rܜ9e0�I�Nm��9�C�,MA��8�N�U9�C!��#/@��)�>[Qy��@T�?�LQ��*�x7��ƈ��uOlA�(<�k���}C�xGT�0��*}��y�B�ns���<����LM����_z�g�N���Ɯ7��7�OOü����[a��������;��dq��]Ft�fS'�EQ��Tѭ��B.�C'��@���~.�ɜ�(+���&�	x7&\�uj}f��J�[��( L�K�Ó��b�v�`�W�ǐW�G���UF�N?>T�U;k=��K��q�U}�#;�a�-���کʻ����g���z��`~D�4�7���[������������_����nr$��[B�J����e��LIn[����&�O��Ni�a�F�9�J��ˉ0�<�M.�lx��	lY���|O�;r�"4'����`}N��](^7�rҼ��i�:����Ɋ\K���Ib�i�L�P��^���x�Rc��W� �a]}�k�_$z�����
Rz�S��~�ב|��� $��˷�MR�-��x߾w�a��x�V�>I;,9��4*�F�]:Z�=���p���or�,d8�I��~��	A?�v��T�D�^lX��T��W�C���\�f��7��4�	z�4ٳ)�4�A��t�B�3��dw�ͳ��~M~�t�9�#�s��0#���nFE�y�����[���}fcy���!������y�D��Ꞟ~c;�;4jG�#R@����}�YLݧ��v��t���H:6_P�"!T>_� ��D��*�V&ݓ�"T���p�!�.ȇ��d6Zaj��H���7��@��Τ5����q���c������g5/z��PZQ�[0;?2e�Ѡ���%x���[�c^:-k�)3[�i��7�c����O��VxS2�,�#U�{.Q,��xfg��JB�a9�T�~�}��_C[�H�T��~�-�8<�1�$�E I����'u�P�d��9��,����A�r��ҕ���^s3�'�`�7XK�a��"�'?�;����7yK���;ء���ֱxe��w�s�l���N�ƴ��m�|�le���BA�i;Ԏ�ck�#��fG#����ƣy�|�|�ڛ�g�V?�DL%�g�# ��?���z�%��(y��T&�:�~ @? 
,,|��GDJ@r�P��ށ�g���u�H���)s�;�)J�ʛbG�ӧ" =7 ��;�lQk�>�W$ �����R��'L�JI���D����&U�>���\�ȿ�Ɠo!��*�,� ��~υ)�LzFv߸�~��9S8�;P�d�*)�ۚ=�>W(~��~܉��C��:�qfV�Ul��(�Z�y���m$�r�6,-�.#�hW�S�r�j�Yj�5,�Z�W<��S���|����7�W9� @Q�P  �X�/�� ��o�� �����x�{g������I��cb�_�b͏�^�J7�n�E	���"��MD����7n!)o�X���!��^z$T��Wk3���<�o�0�,�%(
��k�*IC�M�$���_��vZ� dR�h5���y�hX_�X(�O �7s�����E�U]�����:3?Kr��=�-�_FLx��XSEi2��Y���i|�i�k#~f���R�Z�6c��4l�ܷL�'�7	�M)���ڧsç��P{�����"7o���	C��~G� �X��<�w��w���V�0��<�D�K�� G�&�������mf�����SH0����uHF~I�����7�=J��ݢ&h�D��f(��7�|�g�v��$�&4��5���o��0� M��6��C-��2c��v�G����$t,l&�@0���у�R;*��4�C�[`�kȞ[)ilY���@��� ]��]P����C�*-h1�7�YB��#V�E�)d¨6��Oi~mE
b���k�T�b���?S�Md�g+Dh�頩A��f�:�6�h��!�F��� >L����m�-ﺎ��?q�i}װq��®پ���7@�wPg`���r��B��w}K`��'-�I4~ V<o�,���)�����#�����8�/���jL��+�����8�����`!�Q�|�h����!:����ItW{V��謞f\��2~K�Ry튕�U�B@���N���Fp���5-����0uV�w�@f�"�Ew�`��E��nZ��S�6ɯ:l�/�c3&��KNf��t�ܤh�,�����{�3\�L�\�z .贯�/��+��c��`������ZP�ü�_���00?c��hP?��=wu����_��{f�s���_ġ�lp��Zɇ���t~mX��:���xL� a�[��?{���4�O�SS��mۿ���J���{ͬX�Z5L�����V;�8��������,�g+(�S�bM�B�I^���4\��J�
lQ�~�n��F�;�JDo������?�Ovn!L�sV很\�A~u��N_,�2��HV/�0������x�)c�*���@6���Q�9#����u�J\M���7@U�gU.S�D�����uEqZ:_�a���b��54�
�Vi��k�o����8�b�c�^��4��k����L$Dd^�;;oG$,R�)�e��i�o��g[ �_���0�ˤ�V{��`�LF���z�\��RX��r��N%H�E���;6δ^�12x��q��@Og��\���(�f���m�9�c����]���?�2ݓ@��Zoù�M���2���5���[�k����;�y^�a�vpy ��ߎj��@����������g�V�!0y�w��B^_5�&| z����eT��4�����2#�$> �\�;��<���Ee*��^�/���p�p�s��1o��n�@��/y���h5��uЧ�������h��k�`�z���a�+��]俷���bPh ( �����<���_P��'���?(� qIç.8e��JC)�e������)"u �b<�+�`�]T�g� �)>����w��
 ^�C�z�eY ���)1Jنa^�٣Ӏ�S��� \�ۈ�Ros��дH.;��a�6f,<��<H�WR�k(e���{�9��rv�X0���G�f����/���:�`E���ش�?�q���f��WYv%K�]�T��\F�:M����{l�6��֢RЊ�y6H.K�*��R%z�VF�a'�p~'�xD�9������������,�?�1��)`��:��-�!�$j�u�eP%E~E��^��͂/=�Ar�����KɌ������c����Q,���Ϡ�ay��C�f�^-�r�s��ZF�=�mJ��b���7:/ 5.q}���^"��5\��P��k�	���F�������|Ţ�}2����_�fJ(Ri�U ��#~$�
�Np�mdи���$:�(����`~���H�`\j��3�W���"UO�����#Ek9L�Zr��4L��Q6�ԓ�5K�m���n����C����h鷴A��2/3k�;�����|m"�F1��p�����@Ԗ���&?w�$=\��S�cQ�FJ#��H;��Ly#���T��F6&d��8&e��
nRӴ9I�%Z�N�yb7~Ҵ��Z�f����
@���3�2e���/�p�L-�����i��XI�D3B�N6�f�@� n�f{�w� �E��L��&ޝ�M��&�&	QX��Fk��	�?���9�<�� 4���r�/��fk`s!�	]���2^�	U�Y�c�l���+�y4�oC���^�X��^����Y\�Z�ִ�d-J���{C��5ڙ{�e[��b�e:�Ck�*t��&w��D �o��/o7{4����^D^�+�ڿq�����g�÷5�2	����z�
�$t?H�*k(3��byU�P혗�[�����N��e���������Y�ޯ�קp^�dd���@��#�:��z��͚��h��)��UT��*�o�3$T#Q�YZ͸S9z(5J�ֻP���	'�����5��fK���q����Y��ji��D���8-�@P�^�<rV�9 �F]���6}HFS����?���e	:��(O��1�_ۻoZ>�hC�f	�h�}�U�)�9��?� �����>��(Uf���_k�'z�b@��km%Z}�~~���In6�/߹"�9wb�Q7����T���4��@�Cq(�9�A��z��������'YY��\���ɐ��ł#�5�v��!�\/�o�a ���u����!O,"�����]�Dr#`(�2T���Y��&H5�]Y�v���=��
�j˵NQ2'� �x�P%欉MnRqiCF,����K�8����ֺ�G�L-�Gn�1±�^�>��qjl�r�h+"�����2y�	)'MS1<��ʒ}�%řs
d8��P�/�-L�	�T[,�"��'�ƺ��T%�,Y,�yP�c4�iIA�P^���'nU*:c�/K��p�H�`ا���Ԍ�c_���\ �����:Te'8��.���-�Wr��Ú�p�OӟU��/'�����Ș�L �U<9�~�6.��Mi�hڅc����	�~mt���/xE�?���y6g��yY��]r��]����`�]*�� ��=�0t��bFWd��MU��f]3���I��4h32K�o!���|9��	�}�R����7F�8E�Э�M��޺"���:�e6�k]\���\S�?B��RT-k��C��X	ܚ�6�}5�Z&����Xg d�Ą.aD��XA�θU�1��]������J����
/N�a�a{�wL�5IfL5�>�;G�y^51� 2| t�O.@!0
8'��%�6��b�xa��m�]v���`�r�������ٰ�4��:-�JA
�r�2S��{Y	{�ܹ��p�e��0��0�\������Ǩ���-�l=���5�F�Svy2˼�P�K6��p����c7��I�	�����ѹ�S����^x_���������u-5"��dY_Ĉ�v�������V�r�����W'��ֻ�����!2s�R���c�Xm
4����(x^�~����ےI�>!ؚ���½�~_Y��٠7�X@�̅��y6o`zs�Fj�no���Gm�4?d&�6��g�"����X�j�FMv�$�L@�8�u�&�b�Y7"�]�5�:"�gjH�3�NΖ��.8T��m([u�0����# �((-'C��J�C����pY7�A�	�� ����\�y�&&w<RZ��]�wne�CU�ֻ?�Z�X�^kʼ�f�GI�r�?][��S�,-ڪAYH����ƙ�}�x�`��D\8��\O��m��J�Q���D4}.��`>{nC>]).D�6�`_}!)���˕XM��-=����(y0�J.���^���\#��ю#�zF<��jX�v"��	��>t`�0t1�j�^@92�$�<{'�TT����!3v�-R��rJ�y�|"}Ə\��N2숱����q*�Sƅ���c��=<�J�{�ܻ��?�E�^��]�emRY��yF��]Љ!����B��:ߦ�!U�*�͓}�匴�g`޾�J��M�� ���G	E}�m�C������ϼJ�yB_����ɼ�#����A.�����=c��4C����?��l+�H�9%F�gY�k�Q��3
��ln�s����%�*nm48>�aY"L�:ӆ�.��V�������dc�"�9�zM��t��<��B�{����p��{=(Pd�&�{J_#� ����s�c�$����MT�T�ۧ���L��'�? �(�afh7��E?E�
�p�V꾽�y�B+y�P�"t�dg�@) �qpGG�����I��Z���,yq����f�"[δ�&O�GwJ��E�ٱ/aQ2��W�m���W}}�����{����������$0�Ć� ��"ժ�r��<'��Y�y�'|0��6`��ōܯ��#5����E�t�R'4HR�5RR����a�'�
�OΝ�Ϣ/���[����fw���=y^�9E����w�WO�������$X�:D �c�J�F�a�֍<gr��r���ZE=���8$T�[98�H�Ep�=�����U1��p���փ�U۔:l	^�ا7���X�������fw@ߒf�o��Tb�,����p�4d1���=�h<���G`�ԋ����Ԋ�p�\�˰̇f���йĤZ�3;�f9�_���rϣ�G ��}��O5�����oZ�F�u(�����YEb����Y�"�J���ٳ| �(��!���AKGF�'[,��$	о)\�a�[�t��b#�m��p�bPF���ӘʲӞ��k+�"A)Si�&B����w�*l��47�@gaԁ�tS�\��M�D��kĬb�@/#�aϯp6Y�Qhi�\�ʡ�[  ���g�C�p�R���4����e\�rx�9]������<��7�C�Ab�!oRnn'�}�sm�p���G8z#���*D���$w[/���(a�X�q�~A"���@��]���G�P3D�,{��Rl�������Lǹ��2i�g[S�)U�� 4�z���t�{i2G�n�ҫ\K��I9I@#��=~)��.���G��.�������沄'��.��N_{������U��	yZ����!h�a�t�Fs��6���#-�<�m
�Z�m�<�E�T�>��0�>Bl2�+���9؉�� ն�n@�^
��L�'��-�`����Ⰼ�6eH3�@R�}�g�l�cD���@C{�s<&�ӣ���R�%H��[!����S�E�Jݱ5���
#f��4���ǀ�Q��n��#��G�E�=�d���{!�o��6�M^Z�K�
�W}e�Ú/���:%f��*�c�;��0^S
w�b�AFj�jn�"��Q�8ftQY>r/M1�p`��}	��]�R����@�짢C��̺< �&c�Z��]�� �YV�O�jN��4�](\�b��⸑�����?���h���e��on��s��*�~��
-?%ښ��郢!9&�L�-R'�hF9~�]��?���N�m�
�<A�k?��,�g��m�6 .Q���me��������h���O�'���h��?	��j�1�8��x�v�EIo㫟+^�CXVD��O0ס;b��Bm���o�%�O�&����:�1%����(��U"p l;���6KE�u�beIw�+�*j�ŇP�dA֥dXL���(�䪴d�,2����Ջ!�i[��=f۠d羠�I��$'y�ȡ���3�V��윘�i�XG�o�)&�7��M9���RO��t��ɹ�\دp@c-��O)]c��v
[���tK�|���J���&m�Q�^@�jlѢ��m��n-�[���-I�sa�*Y>B���T���9N܃ܔ���"��ĎɃYa�2�R��7��:�'\U��Tb�:��N)gKQ�R�Mu.�,)�Z�S�R�aE@�t��G9ZF΋6���FO��mk��o��.ʾ��Cc��˽-�*�T�e������;�	�;!�E�\GZ"�M����ړt�4:u���[�q|�?�֕����!I��'3�u���@�o0���Y�� ���7����ֵ�ix���gg�M
Ǵ��T�?5�,�`���B��[����[܄W����J�ѷ�E�5a+��5^7��+�N�$��V�#zC){i2��o<�^yi9+�sϺ��et�Ҿa:{bu�a���|=��%���
�Y	j2i�_&%�.�u����2�Z�~��*ʤ�>�uU�7e��`	M7hZ��t�E��u>��2ƍ�v����J[�ÛZ��lY~<pp9I:aj�h���7O�k���7+�����z�DEq�� �	M�& ,�
���r2J?����~�:�qy����R.S.��o=�<�W�BT�*�	6@v�7��ɭ�q����:h�}n� }#���#{(n����G����U2BM���GlX	�kפ��=�Ո'�,诐�بƄ�˅����G]��6J�mx@�/ǡ��n�i�A]����d=�t`=k�y`B!��eZ��������w���T���V�[�P&'/�-r��#ƀk`�A6�����W5]�`g�y̢�6��6�O�:�v�)�����L@���2��a��N��8��?1�n�̅����52P��K�¹O+���^�2���j~K)�I�AA��)��C���C���ᗗ���B��l�E��QU�0�
�0�M�^D�O��˨g�8�	��-U_(c�A诃�Bܧ:؀mne�d�����&(�IB���n廝�����^����O�+��7��G$p�לɭ
n��Xb4U%40b9����I2���v�I��}#S[�U�+��`?TF�+r�zTDE�?L
�1��h�eY�|,7p��;��o��lU4�(k�8,/*�H��C0�3��`���]u!{ 5�e�"ׁ�����e�RF�����t�b�v���wϊ�)�*=��-XĴ'WKTTb`�6B���I���K�9���,+��:M�t�dS�P�Ijָ�!���>� �K�|T�րZ���� �ɋ�p�̥����+uGl��A����/P�|�NG���"NLD�v��:l}Z��n�}��Ŀ�^��|tH �<��i����EB���=w�ɗ�IA��;_hg9�U��ϜRy��.C�m<pDަa(�$V>(`T��&��A�*]�f����X�HHbS�.�4���
 b
�G+���?�J��S�ɑM0���\W07 �vDAeyj�(U@���4x>�Bal���+�F��$^�F�T:�y�v�o�1V��Z�L��.q�wKE+^{R�X�3�8ۍ��� ���t�*��;|.���e������lE8�1�]_�����l���-�\����D�)���'�t`W` o W��!�#_H�{�� ��E^5�A᚞U|R&��Xۈ��aBi���+�leO�Uby�Z�|�:0�j��P���c��982�0��ˉǜ�H��~�!���M��Y� �{U���;@4�y�%PS{����?}�&|Q�1�w�=�`s8"p\�Ϸ~>_=|��@>,���>-\����1E�/5	���Sa��*|��rk��"��ȗ�x��*�X��@�!<�<Q8PL7/�� �b�_�)+��i*�8,9��(TdA,�W
��9�+�ˏ�J���b�0G�  ���ާ �`%�!GtT��[E�.4d+�l� �V�s�Wd
�S�rn��ZX�{$�K_�^�|����B6(��v�hۺ
YK����}�o/��FP
U�9���g�}���XC�?�*p��ƂZ��83�YJ�v�DT�`_yH�Ϡ���s%�jD\�2��)��_� ��~ �V��U������h��&��Q�k[�{���p�|{��+z���aM8��I-�[/����á�z,�R��l�6����:-ظ��/���6��"���jx>��T�Z��%�[�����Z�V�+X�l՝�>�_�G�IEd����º�%�IBU�0��d4m���5��7a��q��U�����8�jֱW� ��Tl-�P��҆� �#/eH��P��nИ@���Ŷ���i���b�k[@J����[�9��������8j:A��cŊ��F��*�'%	OmMaB�{�t��2����.M�Z��엥��Z�;B���i�����7uz�����rv5C������=�o��
.8Z��v2��:T	vi/��9�Pj���èݠ)9h1� �jl+��uD�g���@�������+� ��~ښ�l�PDhm:}�m�V�p�Y@���ڃ�EJ mP,�}qaw����*���QzW�!I���uR
肅�c�O��V�^����$P�m�Ǿ#�HL�q��${���p/C��� �sk���fYÿ2�:�\9�ru�M�v�xX��JYJ�9�<��V��1���x���+�i9�W&c��:2����*9��[c��c�$�u�2��J�����B�"�]6�~\����T���KK=�A���xW�z��c�_<����J�{26�n�
�o_HA���	��+S�A*����SV��KǴ3��� ��	-@T�� ��9;
fc싉��J���C@@+X�ڢr�2K���S�C9*3�%H�[,fV��D!�<��M� ��@���'X�B��%	B���Z)e�O�U9.hK6���f��Ѥ���n+��*"�"#b&Dtː�B��2;��H�/s��G"�r�Z`�®�0K2����K]n������o���_X,��g��=��QG,CA�Ԥ���j�	���_��͢j}e�[��\K`�/�.�L�P����m�n�ك�T�5�(����6�p]�a�s4�׌`��ayc�
��cW��B��VZ���Jz��{TfJ�3�]�P$�dHY�M�"B��R�wq�c������?gs��4T53.����hNq��8�u@�ЩhD,��a/�h�3���ϣp�\�� ��1/I��`��4e1j�H3tb��0��ul5� h���K7Oѕ�)[ ���j�ħx������.���`�� }�o�ImU��z<O���=n�S��~��X[1�?.�����(�NH�������d�Bڎ�P�(@�U�>���0[fi(��B���=���G�pw�9�����7����>�y.K
E|��bc��V���(��폆sE^I��01�����bd_�+�G��� 5���fg������?����F(
� ��(Xַ��{�5e V���e�̣���o���Z��jw��S}S�%�4*�Rj�9�͋D4=w���f���@�1ֶ�5���)&�1A�_B�&��E���/w�+w�)�`�w$����C�U��a��330�ԼD�ip+G-�T���e��U�{��:p���'(l|�e�f�x�@�Y̖�wXA����~`��G9K��T��9�!��K�K�J�J�Պ�W+#\bVh�� �y�_^�-�ŭ~f>Ōx���q�K��*PbڸSx��y �s||��6/��<�\E#�������L�鈭�h�]z���/��XN��4�[�Gެ���,ۑ�\/ &�Is�'�UhV+��f[�l�`��^�>���ͼ�O�pq�ԯ�Giz�GHȒ|ȋ3d�
��Qؖj"�]R%���2mM�}�+V�@0��qX�c:˷}�@Ƒ�Z���A��TV--3Us2`���XZ����F|���N H�b=�L�S?(A|�$K 0�"�Ȱ��"]�{�\�[���:��U1Ø������SD��ldb�%�����������?	���_���lĳi�H�,�h�-_ݎ;�"�=���B�X���nD5(y#_k�-��؇~d���>z���X`�;3�Ag�U��z|4;-6�#��f��T��#�@4���B��\a�-K���>a�x5�Y�(��p�'�K�o٣�Z^}��OlZsHk�(0�V#�j�\h$l�#�3A@N�1U���x�mZdi�\��F�]���!|�y!����f������O�|"�+W�Xh]P�(|*��]������[��y�-w7���� �D|��B�}7	D���B+>DE��dks�$м��ʹ}�"UT+]����89R^�P�d�P/�_�d��*LU��*��)G�`��h��ƚ��J���m� �p���e��o�K���|���Rt<>LJ�I����,8{��<a�fd�Q���b��T8�� �A\�p J������Cm.�,
��z|�%�*_�,�"%g����U��Pm�)�+CXAKa������.m@@U*π�,�0�WθƏ4E�#�pJ���E�۩J��hm�a�A������D���F�Bė�[��/3����B��,K�_0oN��=GA���DqF��߈����R��D�bUF�	��Xb��,���l�-�;�Sk݈�T ��'�P�FO����E�����G����������T���N �^���P/9�B}�x�Ehm��9�6d�%Ef
�j�ݷ�Y���]B�`D8� ����@���@��o��2p����(� c!@��������UM�"kSY.���7Sڏ ����5ڂ��B �)p�X����������ەFM�(ܳ�����oU7�
䮵�-��6��\U�Z�0b�@3���+�oP5e��1�,GP�hL���|�L�$R���"�ʇ	w��b�
0��(4�6Z^N��]�%��&���͜@�ZҼ
��#�,! e��������d8�-6'�1��k<���f��f�r��Oc�:>P��'�#����`��2��O?�)� i��4��U��<��c6�D�.  ֮T��DIyU�E��F�����h�`���\�[w�VQɀ[}�Ql�v/� �bef�p85[~q������ί�����[����c ���(j�w�B���vI�y��qiC�	G�:��:�X$!�PE�v �@*,��"� -��|��r*r�"�vE�5hm�@���~Q��!b&�,� �M�����ɒ��6@��sw����ur�&���1t%~A��|�Un�?0����.�i��K)۸,���"jf�8�Y���q��RǞdlt"&}ܬ�ޭ��4X��˚g��HER���+J��`-n%bU�m�fl�nB��*���T�a�������̿�k�h�,�ڱ�����=�h���(������G ��=�j�2�ܚ��EF���gB�אb������K��w�@H�T�81���XYIi��p�2F4\4UN�RO�ͳ�`B���� N%��
��]/�g�W	��˧�Z�_1�9N{A��SޣuG�H����,*�Gm�oS4b�j�{@��fI�ҵ��o����4F��<t��� p�	m�*�%�A�_R1�0�|�Pm ���' <�h��c�V�˽=ݡ�Qb�YVr72��� c+[�� Q���rg�X���+��r��ze�_t�����;�(�db9�A�@��h�W� ��١�+ZI�C�+`P��2���&Y���k�J�Gז8��F��7�ށ��}�����w��k0k�zLK,U���Xo����r�ؗq-]�
.1� p�0�
�L�)����R� 9�[;���8���ƭ��4�8J�FZ@|����Ӊs��j6W�
������d�{6�0��o���@��R;tBsi2�ۉ�B)J�X8�{��j(|��
a�³w���% �v O<,����I���ZƕD�v�����/R�S1�/��ێ��+u0L����<�5MT��ZU�]�⥮z%n��ʈ� �f�.��ol�F�d��-"]����`�`�Æ:��@]���+,���a���eb��s]ř)>?� ^�TN�r:�K�NQ�XT�a�[ �*���t"	��@���v`���P��P�av���L��i.�mΝ��H���hE�Pڲ����Y�n)K,Y4V)J��k�}R�,�#@� �Y��*�Is0��(�Q�%w���1�:���AΚ���!ܪ;�<���4w1�ٹ�ލD�6��y�߈��[T��5�:۲�~"��>h��2����F�3���U�B��𔂫���r�ˬ,`���x/�����Fʁ��j���EY4Pp�BH�h{�e�$�'q��w���8�!��A����L��\�D\�m)��nϑ0�_(�H�ep@�}�@;���t�2�i@�%�Tʢ�SE��0#��l�6��+���vɀ�n*=����j*���-�i�{�}EKD�����%�L��y�5E��(�|��m��@� w`��ݔ �x�� 'ɕA�*C�#S�>���w�`!BM��y�wM���bQ�aL�������9 �4{�\�%�,G �ʬ�cx>J X�ٚ�0��S��q�%|8֡�g�Tg�X���T#PhX3(�����m��.V1��*(�AV�'����O�)��k�i{,��Z����2�WrS��)� �2*��	���2��
�ɰ�:��*� �'� � :���C�����Ъ���P�)Z���bл�E��=�FP�͏A`U�]���R �������������
Z�1��<�������BT4�<�x�W���6:�=�6��|;4^/���!�j��� �P�r���R�#g!<���A�#(L?f^����5�``�6O;�m?i��N�K�/�*���Z�"��9��?&�g��_�����.�*��1~A"��E΢�\��NY��_/�K1c_��J�Sߥ�5 �I�DF;,����*�	� �*��Q�G-Cj�$"ԁ),	gf����
ٻ�Dʿ�Ç�����a+E�,��r	Z��ew?��/�bgA��F�* ;JE�5��ju��Oܗa]|	�f�̷���ؖ�����Mg1o+�/{�N�9��r��>s��F@������@G%�֥t����|䜔_�J���*�
��Rڵ/h]����,��O��~��{��fظS��ʱg����%�X�hl͆
K;UNJG�V�Z�3���m.;�\�;�݁^�+�ƀBu`�G���P�%�D��v���e����CA|��/LfŹy̧�c��`��7�3�C;Ұx]�� 0d2:��H��Yy���Z�❌WW��J�����&��-�����W��+ga������oo1H�t�3��8W
�$*v��� p��+A�.k慵FMc�@
_7��#�7dm�r�-�T��ƾ�- 2���� R�n&��
�%V�!��r��v����r�H0uo�@dA��6k�Gi+P�?yp� Z`�;Юb��0x�NR���qpS;
�����yo!J=�b�U�܂��@cȘFx�arO7{;A�=��B���<@/☭duM4���N�����1�ĝ㈞B�Z��ҧ��w��,Q�ᒝ���}��ߙy�D �f��3t���@F�E��yH��k�;+�JY�"F�
�'z�r6�J<�:0�@�Z�������8�,$�kr��+O�{ѥ����"���e��j������1��$�֪o)w���h
�H��1T��OhD���q�
����x��HL�@x�4d-�aXNbօ��|�MWL�� �����(g_8k�k��L@��g�.2Gc��Tɖ6�<��t4SM���=��C������� if�1/���ڈ�J6m�	�J���8�9K�ʰS��_�B�ħJ�h�_�4/��k�sd�u|�B��b���Y�`� ���MޒU���B�[�(~��5Fp�3�|��ǝ�5DJ�_���2T�~�SDr9��,K�^ �|؉�%3`����Dd:�=�

�2��2����[�ۍ��%䡭����pX��V�T->q9����-�
����]+).ep!��U���9���qɖ<Ѳ��Xm�FZ�(�)zT#b�{�j�P4¼�i�k4C�PG
�30L<Q/�mE��
q�QOM;��	2�恈3�i.%�P�=_m��d��Α�NK�F�0d�s������KU d1�C�<,�#OeTGK�B���5b�J���B�{~ �2�щs_�+k���m������l�(���pL�Twsz�Y�b�k5����4�V�+���d��,��	���-g�F������ݧ̫%0u�e����I���v�1���q��$��R�V%�C��m�v �,i����7W��&�%@������-Q*��*���Su[�
��i�,�U�QW�lHY,c.h�_{���C�	��x�Cp� 4�su���pn؄mm¿�KGuG"��܃H������Ԋ������R�NNЮ>Di���7��CȌ�Sd�s�c7~�1)h��.S	�*�\��J��Y�R��p� ﹋ �vG����������� �YH������*b��Ep;A\Ðo�n(o����e;�r�fL�����n��� s���wQi�V���|��cj2 i6w��!�ª�J�#�n��p�� GI��� �"�~#�$Z
X(H�m�X)Fj�/�o����=�ưv���9���@L��v�/�y�l(�ڕ����<�c����x��D��7!��"Q�e���D�IE>�!���io�� j#P^�{�l�@�G���#��y�d���b�`������J=��)��a�I��f-�<�v��*��*w9���C%�����uA��x���%�|EK�����k�T�	I '9!�A[�,@��n�K0�3�B�Ç���g*ƿ{x�i��i�6,p�T�2�^��t����eyOv��9X��Nb\�v���|�D�ʫ�9�hͩ�����qU|���Kk,�I�)�!����E`=����x�J�o�/�/MQ_��y��?�:�Qk�1Wp�"�k5S�W9����b���.�$:E�'��Q����p:Ŷ�L�b���_"03�%�a��i���p�O~���T� ����-�'�8��b ���1��;&&�kو�))�,��H7��ut7�X�1p����@v��:/���� ��a�	!��;p�l�x�Q{�M�ݭ�~_y+꽦����{�b�|ˁ`���I�^�c�p��.�
T�JVox?�w�ݬ�ޝR� ��q�̓��L������u*���}�9�x��ġi��y��H�ߴY������'�����Ccz���,f�W��M�#�KO�� hA�~��k�39+�(���Jj\X� B0���G�n6ogEJ�C�(�k����4w�J#G�N3*���c�+�"$�G�Ut�����wTVf�M�q��u�J��Uwv�#��5!��%_�\��yMsm?J��P�#��n���A�	�<�s�b�L��� �8�4Z9{J�j�,�K'�@���,�
@&)t�_��¥�Ik�|E�}c��_�X�����l�sW==�d�j�����[�T�\�V�{�V���}��ʀP�����7NP!^��V^0��Q�0���k`� ��|O�O�Y��q��|_�� Le4�*���t��Z^�am�e�@\��g��F�tf�2k��.�^;{��+oi.[�S�\u�|�=�����H�����Յ�y5W�]z��kp�ͪ~�Q DLW<�|�@�O���H�jm�Q�-�;2w(�OA\��z��]��1�}߆�� 8ӫ0��3qDwm}�0�������5+5� g^�5Qqľ��֥�s,6�@ف�*�b�.��ܨo��\�Y�s3�0ķ3��(q����o����a�nx!��?,�����	N�'�j�)`w���Nq��t�����@�6�D-���@;%��k�V���@����C�n�PM�3jc�c�R�k3��ƺ��,�_1N�֚��E�,�$Xl��y�g�/7���o;�����4ȕ�����J�r�kS��0U���0P�'���`C� ��*H, ��	b���d�������-QV΄��/%�����G9����f��W8��Ȁ�#��0�S�, q��	XD�c"�ʸ#���T��s>r��k��� �������ܤk��Ls1� �o7��So�X��rJOx�҇2�1q.|�f-^�I��E�LF��r�g�o�YR�~~���D&�������B=K�\�f;�	����E�``�`� ��U���m/��!4HR&o�6�6�L�(�&xD� �cq�?��	�~a�r���.a��	��4��C?X<ee�:)0ٻ�e�C� �ҍ���T ��g���i�b�}V�Wk���P]}ng���ǅ�j�i�^����
�~���r�|�97(�>�e���sP-�A�ʺ�k�q�+��j֥�D�7�+�MC}�b��'�� ��j��a�1��A��ɍ(�#��Ζ70���7/5/0���W�Rԯ�&z4N�QP�K�y��.���q�� ��7|�� 9�v�2��Vb��w��Vɕl������K��D��%ؗ���S@�h`0�M	|�t]G�g�¤�r�:A�Ѳ�0%w
(�������-�=��"*=�����j�$��1!Ơ�ul
F����{L���Y�Xb/�:x?�F��&�z��9΍�."�>s���<��K� �ə�ʽL��AC��q�����W�3�(�(�xZ|�5{e^��p������WxE\f<�#�1"�y"���
_8� ��U�913J/�Ǻ>�\Po;��gӷ���
�Yema҇����w��S�-�V۟x�����+�Gʉr��A;�1-G�]B�B����@a3�?iQ�l���n�Dh�a��u/Q�B��D��rn�����[v���� �?i%�j�F��8��KX#ىw��֘��Y�r�on�s��k\Ą]>Ő��U,^�s�u�~f*-nb�ln�4�L/�eA�M|ÈYޢԏ�E��w��,.�G4R}�)�O6U����^p91������"W7���.]t㶢_u�����Qʬ�Z�N��*���kp1Z�\7,@�|����6!G�����r����//�#L��f !昐�5y���[�+��=��O��s���N�̬�`pe:{�򁥴�0p��`�{��xb���r���V��p��-�j�`Z��qJr�T��+˼�8��Ҍ��6R{tS����g���e��� �s��Hr0��?,¯�W�wÔ�4��݁�e�f�����W��08�Ȱ3��D˷<�b�g��=���,OΑ�:�3@���b�B��j��1*�e�Xy������з��kV�6���ģ���2L 	�nV�؉p �F�Sm���������M�BTl��r�2��P8͈�+��� ���
+r��x�H��,�W�}c��cE�et@��+)��
Hh�p�0Q"樰B���y�Q?x���?Y�;o$M�S�#����k��3�%-�Jw-�PKkd������&>�Q�)l+��U�{?��衜s!�+]��*
h�^\����XW�1A*��e�!}� a��Q ���@7G[�&m�S��Z�*��V2��}�d�r���9B��P ��G���R��,��9�=�NW�t��_��|�6�3Z���R��#�@�p,0","�[�9�����B�ಠ�@��� i���� Tv,�q���}����75�zX�A�H��AX�8��T������QsTAb6��7T�%(s$�@b�U$�x' �-��)��T�ƭJ�e�\��J,������e�lD+3�c� P�����w���5��K�kdc�+Z.�[�s�$1�h�KJhp#w���/wD�R�&aQ�G�#,PZp%)h��.[���d��G�S��/�] �PR=�c )�e�X|����	�� C�J�
�Uky)nNC��"�atА�1�j
Q�z�{�U�W�)��1�0�Q��!u6n�*�q-}�Lc�����c*���jbU���5~b�aĨ=�Rqa�H�b��^E��%*i���j+!]� �=�Se.�+X��˹���[��2!���LJ�i��(��l��]�8D}�Z�zxE{g�_�Z�����-�X$�/&�q6�Ɩ(�T@#��������x�x�SBr��(*5d+��ۖ�P�!ZC$���[�xj2�8+p�9<v�������Q���蛨)أWKuiR��5߼�j��@����,�֊.��[c���e�F#�6h�V�ۍP��Վ!i�ǹ�S��,��O�;� 'e0����Dn�^0�ZQa rE�-�W��� �S�|��U Uh��\�M����B���X����U��Z�E�D���  �3vLup�3�nsɜɧ;�@�M�����iv���3s����a(��R�ۊ@�*�;1I�cb<�1i��ıO���1����3:�%�O��W.M�Ű-����hN��yn=ߴ;�-~P"Eh ��J(��GI�iF�q�nP}z E�0$z���� jQ]�<`��*��J%\��11.5��Sw��3�K"�����<����S�Huꌅ�ۘР�d�
g+X`�/i@Or!6���:�����_�A���F���8f�&��@
�Lf�0�\^����;\yU��FF�ɫ�W�P�]��x
&�7,Ca{�������Y)oѹ���e�$�Z3,�@|�Ƞ9B�|�)�HcF��d�Kn�!�Y��2���Q�~��S�zZ�Y;��y=���ѩb��c�eh��U������f�B^�z��GyCMlR�y�����͝���ԩM�>�����p\�(N��Yp�V�M@.���GP�r��F��4�s�m��dඏ
����-,����T)���@�U:˪&&���9�e�G��ь�4�'	��`�f�I����j���Z�4�w��K����j�6_[�sm��X��4wMb��wU8ϼ�I��<�P@�i|�0��2��t�a��z������b	LC8�[0�]q�a�lЄ�!g��Z-HdG�4�.�k �EǸ/�Kj�ɬ����P_6�D�C���XJYR�)Q��:������e$A;�$Op3�M��,v3Y�MH�����(f8;��Ȭ���n#�(�Thi��U�ƍڻ��P$�ԝ�<CNG@���+�ZD+C��zS:�)~~io]�,���/Ty��9�A(���������T���q8`��k-FѝEԹ�J��g�<ñ@٥�3��L�(6����)��G �z�oD�>@/�\Ci_>;+�Ӎ9u\�-%6F���%gw��Y&5�H�x
j��Q�n�,��G�?�� Pb�������d(�����2��E"����H梛��y��T� L�B��inŠ�%�B�}~��鐴��̲�)oV\�5����^j4�T12q\��3����3�m$�Mmor��ww�&L�!3E�[a �Vp��#;���w���� �V's�͖��=��b6*��#ml�Ƴ�]36G��2��b@
j�b�P�"�uz�1�`ı��P����}
1�d���Aє�ʄ��B��B��(�ņ��T�n��Ar<�h��,�v �Mf�qj�G�y?���>�K߳��0?��լ5䆬�?�22���=��+�ޛ�lCR�����wR�Yc~ǈ��V�#J���J�[�C�Q{PB��70���#H��W�J$o�3WY"����(�Zi�	�1��R��I��X���� ��J��5]��S�>q�S�˗틺��QF��W��
��_�k2��T J��o7q��:�2�%��\���	��E���<���_�)��@)7��g�	���`qU��Y�����z���*�E\t��I���$�U�;�h�re2�7&��r���?��1�2�C_�hGu�hjo艔�,�XC�wPSm�GA���&*����@����))��R�x��\�� y"=��@6����-YE�� ��ٳ���\�v>҄�Z����3�p�6(�-��5�Y3P6[�y��7Z��%� 1�$^�.~��� B��e�2wC����W@.�i�h�Y.-(�Mܤj:�3���ڢ�\Y+O|�*�����R�X�,/h�-���e��j9*8J���4���8eX�?K`k%�ڭ{�	(dU���7v<�����@�~����?���� 4�UO�����t]�JB��O�?�W�e)�V��ST���
���:;�+ *��sKx�X���o,4���U��-��@��@���٧_f�O �9����>cu�b����
��� ���� ?� �5���*T�R�y�9�p�5��J�*S	L�S)������ʔ��̯2��^e��K������fffff{��+�Q�p��|ݱ�S���@�rsс]z��-4@�F$��a��f3<]��.a�����Ir�r�b1�*T�Wܤ�{JJ=��+�S��;C�u�N��$��\`""�j*�.\Yl����oB�(t�B�0�j%����J������W�X�X��2F���
�+�R�����$�F,�eH3H�7(��jW�?0 xA�sp�*&,Y�VWJ�c��(Uf�%A���*���=9�n�o��A�s��]*T�R�T�]*T����X�Nw��\w��2��u�j�Tu�㾗3�_�.P���R������S�"��v��K��0��;��pJ�W���N�"KYK�(�T\���Ï��WC�8#��oh�>;Y�l��fWR�KR���WE�����R�:�i���	K��%�OC�jFdw��u=�讕�tCC�G�ipW�A�����(ܶ��fz��0�_�?Cu�=��>�芔�xo�Vv����)s-q��p�PR���w�ҿ�~%�R0�*n!]��X��/�/�}	}/��/�|GbX%��M��[{���;_C��3�<=57��-�T�]OYҙL�g�˗.\�r�ë��t��C���+-�.�d�d�K�.\�q�nǢ���"*����D���iR���7�[�r���\�r�\-�"�BBsӨ�؋3���Sq<�Q.`e����W��"ڳ�� ��Y����x�o�����[��zOMB1�G�'Kt�,Q-Э󝣯�)&Շ�^(I0��b�<ĭ�b�B�/0��=B����gW�'FTow�dwR�sz�y���P���WJ�P�/��貢�����:h���w�P5P�F<�c��۠�����15-9�d1���.��}&0:��<O�7#��܆"Y�tz����Tw3�PE�E��g0�7����x�:}�Y�WE&�-��= ��
�]���$P�u2���]���>�O�����$TsH�l�T�ۥ���*㹼���Q�:�Р���1��������8ugfzif������I4J�r���ӲkAR�]x�X�
DN8���*��l�0u=�Uˋ2�~�߭럺!fT.tQ�p��6�r�^�m@�Zp�D�10�'��gw���zo.��jT�_f��R�J��d�R�~��I��6?F�T��.\��˗�~��뢽�J�����_ᄾ�7�;�����z�Z?�L�O��=$K�}_���q-�.�FB�r�J�Cq��VA1�G�-��øC�Sic��nS*0�_E���@�̸���Dj�n�eLx��HC�t��LX1g��0 ���Q��&="]#���tW��ۣ�l�Suq-e��>�],�0��5��HԲ�La9tuC�&�+R쏣r��G0��u~��֥tW��C��Rӂ(�4����Hܻ>�����������T���Tm*Z��� ������z_K�J�+�=<}WJ��~���F=�Z'J�w�{�m�i}��~��EKM_ѹ~�+�[�+}._B���:_��3?�
��Tz'��*WE�z�nC�_F/�]���\[/�����X�Af���j�?xC�D�E�^}7ӿ�z?�Ќd:9�So@����tq�D1�+��;b��{�N���6�E��4��EK�E�---�il�Z[3��P�ALP�euz$7�5�ܸ�Ash��Tl�Q�e�P��Ńg�ut���F �r�1��a�5�,����./����ҙi]X-��ںԤ7ѕ*WGR�@���32��AKKKe�ٙ���o~�l.*s��ε*W�����XS��[��r�\ t����|7r�\Rάo��w���zs,���(�RRTrM~�����(�P꒪��>���>�2��nbf�m0o���Z�B��K����z��4�lN�<?�:�?�R�\��KE��k��_�=9�W��ܴ:U��gA���?F�U�C�*\���%@��~�:���=9��� X����Ố�ˉ'B,q ������_�@�k5�n�:2͗Q�h��X�����tz�9�r\���~�:�ι�s�4�*�~���[��Q"�%��Y��7���1%ve9���/����tQPw���5�U�f�tz�����X�v`b�z�]�%����u�5�V�z�P��9�Fr��{C�ޜ� H��V��
t�k�O(�n3Id�%�QK���J�搎=<�tzߠ�	R�uYr�O��D�WP����4�5�a���1xz[Y#��F$���������[/�z�4�>�N��)�G�tsl�P�-�5��Bg�1�ߡ�*Oҹu(3�5��Q f�ԠQ��^W0�$=*RT���(�-�33�ffffffZS)���KKJb���G��M��f����^<��z��%zGEJ%J�֎�ҥu~!ԇ��+�dM�2��Z��J�}C��\����S����uL�R��^�q�}It2�E�yT����p�Ȕ�0�0T�\��$��45�������EE��m�� (䔥�I)��l+@ŗQ���r:�3��q$�{�޽��]�]�����޿~�VU��#�I"<i,]�����׬�A�ф3+��=n!-i���ӹ?o��ȿJ�ݬ�K�t�,�B�(��`���25�to���7�2������f������e�dfG$��ҫ����.��;v�_�����/�ɺ��J��t��@����0��/�J�����hiq���q+[��!��x���Y�Y��J��A�77�R O����z*��Q�'t,�8�XA�^���ML��<�+qA:���|<�C�����K����O5���u[�^~�>F�Kfd�$u�T�`%Ŵ\GC �씑�'"��/��s��B{��i���5#( )�]����$�c�|�g���]�2Ѝj�j�˱%�S_�9Cu���O
.���YΨD��/1+�(���ong��o�B���Z6q� �U!��	<���Qp��W��S�==}��터m��Ùm�V�Kފ����T�.�E�m���	6�Ɋ��2U
W���G�w����vVџ+�T_���L��%@���Չ(�5����:V�*^v 1�VP�ï�q*���K��q����֚�se�(�� �\�ݽ�^�_^�ibj�ς��� Y�p��)����8�z:֬��� �J���N5����Xz\�(7d���Q�-{��w���)r�ɶ�J7�PG�� ׀�I'��:+5/�������X�����]3���O7�cԬ�����n�y�����$m�Düv�Q�)�R�R{�jQ��T���&�;�[�d�]�戠���k�"��Fo�W�f�I����/SK2iɅ
��ن�>.�N��d�5���q_���Fp��Y�5g5֤n�[�Mx��=HO��Hi���K%f�w�z]��x��V�(�Q�/I{"(>�B�O%�FcP��!���9ON���u��*ͧ>��#�X e�]��S$x��N0E��&Cףm_��ӝR���-�^�t�@�9�^���;���O��7��}�8գ�+`kFa�����y�"�8�!̩¬śc��"쩠{�RS���x,q�[�#��)��_��C<Z�w�T���P��&q/�X��I���V����(�ʙ@2A�jI3q�T3��.�S�(m~�_��b./�m@`����X��Q����z��όa2��-���� ���l�"G�����)(*f�[yj�tz��B�+�RP��-p�����bq��gN�_ߑ���Ȩ��wÚ��y�L�?`#�tF��B>�󗳳����fh�S�|����d����]�W&���b@ W��_�c���(�Qa�v��SBVt0z��w�;��L�@r�:�䃎H��8H�C��ԦQ���ֻ�`5d��x�tU�����7�l�5Ѱ;�ya��e�*/s��a���	\	8�ĩ�p��������������)�wǓ
<<���6xb ]ǔ�Z���jw�%�+��4�i�¶h��������Ga�wTvu�krf�D��������|���ך�9!>;�"&yq�f��65�D�t�(��5ܯ��[.�jKu��������E(-�.�����h���C#6a��R�"�B�zhT)���͉�y�/^�����E�Ӆ(*m����W��>��n���"��lh��D>NH3\F����ku��f�YQ�|��H�Bp[3��%��f�l�x8�#�7ԅ�?���Xc�-s�dyꃒ��&�WSI�$�U�a~~�DQE� �m�ڟ�=�Ѧw��Y�"�����q��������&�0[��Y�he�v���������6�������`���@}p�n� B���Yf�Mo��\|}V�Br:/���x��Am(�c���ޒ�S)mk�!�
�}�� !����v1�3��=���}����#@~��������;��S�x���ή��bqP-͒!���U�/�x�<�!G�@�A���W�oӶy���y\z��}��q�p�W= ��b�/2��<5W���"��խ�����抮�4��
��U����I��A���~���<;ւ,�*U�7�m�|�#V����� Y����>J"�G���\���F�p���2]�t)"m���t���t����L9?{<�Ô�p�4Np�v�����#�~�É'��Jߓ�P�f���iԮs	��͍w���L%�SFѤqF�*_��z���7�PK   &��T��beY  �[  /   images/c5cf112c-a0c7-416d-8826-4525095e4ef3.png�{sxeϲ�m[�db۶m�v2�Ķm�ؘ��ۚ�����{�{﾿����^�wU5��zuW������6 YZ\J �hAh��w ���������)����������%�����������-�7==#=���0��:@ 						��������������K@N��G���ILKLFAIEM�CD�H����+�׿��@AA�Bâ�¢}������>�(�A������|�  P�O	�	��`P� ПT�O��M���}J��������:��
#��P?�" H��~P?�*�A���  ʨ����S���;�����;�?�wH��1C5)�4y�䄥�����+6�d��Jh+��  h�ȑ]���E	M�� HF��Vϊޗ.�B���ֈ���t"�!�����,�,C��G����ݹ���X	�>o�r�� Ҫ:�Jc���)��k:��O��d���H��ўqG�^0�+w}�Y3�W�z=j�v��������~��z�_�*~2�2t�_Cy�G��p�P$��fU&k,��7�#�h�����uUd��5i2����r���? �A~O>�_�d��s�a� <�Z�ݕ;�4O՛�5���m&�,rD�\b�k�_�qWRn�H[�c��/"�vn���'� )�  ��z�iS3:��:��~[&�7߻���!'5W��-p�G�G��K��NVO���g��]z@Z����a�H#/�;�5�uYv�㞸D󢥕�q��h�kًV��k#�m� )�V��H�[�}9�L��;e9p������ �@4`/���v���|v�)Lip2!�tF��(�˯�L�\��������U��7)u]��{�m��}�H�����������'N�)��j9׈�>�ʵC�0�*�ф܂�Om��׋E'@�� �M��\+@y���QȚ�0#}����#�=`Kִ�B�)�`5������L&g�����)��up����r(�mS���~�e�M��sNW�<��x*��N���,:"�8\��~���r]S�q�mj�f�+��7�'����F��j�5�t�D�����y���GIԾ�n�leC5e+@�j������I�do��M����H棍M�	��ւ���I�K���k9]6�Z�c(�d���k������Vٻ��e��dn�� ��'��Z�<��N��R�\�?*j ��l��ȯkP�7�a~f�X��������@Mט�Qʑ��YOd�>�ۦ0�j���Q�e��D��˛Ջq~ �B2�R�Zz:l��,�4\z�?gQ�����:�txg�����Cɡ��m"��R&������!�q�
3�7C�4�^�r��/�5�^�����	�O�!��&o��`�~�Ύ��eG��/�^��9�?H曕_86r)�c��t���Yʚ6�����cm�^ׯ�ʏ����f?g��W�i���{SN�l�3}�1p�~����T=S�����W�^�J�Bo LE���w���M*�!6�詗�����x{�T8���w� ~��r�-���1���\�RA�
yy�`;~�hDo��I(��q���~��	"
���7��z+��r��G�ԱYXbP)��·3�{O�r_��Jy���2߳�EG�B�Fk`��޻�ցt��80�s��FH9T�ˋ����Y9��}6����a�9l�Yڒ޻����v�n1{q�b����?��S;���~Q�=o9�7���?I�yD��e����ͯU��sN(�a�M�/�E7^���-:�?;��-� ��V!9�bg9fԚ�,�ƏrY~n��[��;�yv�^6������U�����*����jչ�\.�՞�L��o�J�6�$�8fT�dR��"��]W,t�_s�:3��m<[l����B�=�t44
��p&{�����g�=���9��֠� �����w��X
��J3*��rE�Ǥ�?y���M!������eM Kt�my~�>==s��-x�e؟��]?}�͒�z�3��x�U4K�:��'���n\����3do��[Z�;.�1�^\�nW�.kM�L��F��oo��? �����'�l*�u��0|�f��ʓ��:j���-�Ւ�=���v|�`G����0(�5ڭ���)FZ�zx:����h���  �Kc��E��h���$���
~�$�&�S!�-|Y�[���������ƠG�����!���eK|Z� T4tFdR&fH2V!�/l���g!��lq!K�?����k��B߃�'-gb�����/�R�ȣ����_%�ATM/Y��x܅��V�BQx���d�7�M��f�"��b�%��I/pb����i�b�ay|࠼�@�����q4�� �d,�H[F1��~��fm�1���v���6q	�uC�W;+�F��{��z�:�(R�g}Ćl����_�!pC��^��/�T:��%P�٣����Ub�z�pY����3��#��F�BW��#��l5Z��;���>e��s~֛[ZlzFDŗ�m�X���e�긙H.��bG�X�B��{D�}�ƒ���T8>s�c��>���9\X��h�ܲP� ��c����D����JhiY���)[T1�LvqL��+-VQ+�} d���LRNN���9�����u[��n����elI����f
t[hک��9,�?�R������t"| 2�i�j�����i1���$NR���olѴ��v�������Uߗ�����u�nX�~�ƙ�����������x�ʶjSCj�<�[����-A7�H��ֶ�n�l6��C� �5ڵQ��4�����aY�]G�e)ۉ�g���sZP�g�퓗 ��m�W~�Z�$ց��ܧ�	;Y�� ��Q��@S��6��H��=md�K�������tS�rO�=��d��,��������|�L`����/G+G�t�(����>���{���`��³/.���p�_/��V�>s��#g���3z��ԖӦ*$e��_�/ߕq�NrZp���O����-�z�l�@�Z�/�N�dV��
�N����ɝ�O���G�#_�A�`	K<����dxJCV��7HE3���P�'���&�G�ͦPB6�U�:�?���^��F���ŭ$9��r)Ht�W�{&�K�8�4��ceV�׶���BA��ה����ġ��	�:� k&��T
�lftgx�9s�^D���,�
������!��]N#�a���I� 5����-%D�a(Z�5g�kwj����?X���0\ �TY�:�>�'�t�����9-]�_�VBa���'h~$r	�:(�����X�D��s�N\�:��Pe�@�r�����םb��Gc��ZyQ��(E�;4VƇ�6.�3+�����V9{���Vt��<�-K�K���G�Y2��E��3��h�G���o���k��p���4VC�%�ꊗ��)�����C�7W[]���"��7u,W��2�����0˖-�\��'[�h�_�ȫ!Nl@���Y]*���>P��s��t�p��T^D���l$�XG	ڡ��7���{t#�?��Zֱ���6�9O�Oֲg����| ��%��T̈́�d����&�d�d�uE�#��|�9-���|�;�wqH�BG�$Q�? ��&{��d�>�$�#=��g0�`
T\յ�A��Z��{i�$摯4���\1�#s;���<}�R_�iDj�um�[N��S�l�M���&]�L�����"�L����MB%t}�/��%Be��"C�!��ϼ8/�_��Zs����d��!L���X&O�

`h|����5�32Ay��]����3*y6�?.$U
)+5�vW�C�Sq�ל��`��X=w-{�kB���K�I��xM����uJ��~9�*�8U���}�/�%?�������4W��D���C�����.G���P�2mbELX�BKX��#�'6���뉁&���O�>�{v�T����C��e	�*U�H�s�նx�wS�b��*����D������w�x׎�f�S�Y0e;�e=Dlx���y�)rlh���w��d���\5�4��Rl�v�t�L�7Rd��.4�"�C�����]�S3� �;Bl�lc��"?��;Z���Vq�D����0�N��o!��o&ǭ��'��eB3_>��9q��0�d��,���T �[٧�� ���/;��Tp&d4Ff!%#tRbec�@a2�z��l�Ϣ  #U�K ���%���ǧj��>OUP�?�:�Q�3y^�,�utyhĞ�y�h������s�?|��JG�H�M-�Z��Z�r�هnN(�U��fU�0X�4��W|T�N��Z6�eK�Fey9;�|�c�\�z��a�(X��0Yb�"�h!���ѹ�]ٔ^l4�EU���9v f0�	s�/�{�:.���i9�� ��6!�e�yA#��5���3�{�Xڭ@r�
�SaX?�Z���!(�I��u}׎D�� �._��Qs��>�-�x:������&ɜeN��v�u=�$�6႞�7�_�$l�3��e�8D�*M�[E�U,o#�85G0G�5P[c/��R
)��(��^D��i��V�� G95��OU�]�-_��[��~!$\+��+G�س*��?�'D@��ر~�تCL��Q�n����[��Y��m
��|E,�ea�Tuh�2X�%U=TS|�m�8����4�ѸJ2�17�KE=I;�>>�JM<FV�{1E[�����'���Ďu�A���!BW�=q_�s�s�����/m�yA��ƍ���״͉H�~[%.
���@�,�s�1�1��������~�z��I(8�&`�Uj.D�X����Y�~}��Im��G_2ɝM�"Rb�U��~�8i��"1$,�7�EM}y�}*y�Z:6��őL�w�D�d7%�U<mU�����T��+��b�Vn��n���E���ۻ�x���5G��J���4���b[&�ixQE�Pˉ6�i~=�eS؟��C�:֎(���[\��3��)ȥ��֊K1�[4�mX�[Lt=D=6�P��X/��R\@�R�[�<���h�;(��`g����1K+�gHeM����z�0tq�����-��'̧�C���ǩY����R�8g]w!��@�F�V(M�a�DB/~�J�B����3���Lu���8�E��o	�4����.�P\:���v�Ao_�r��kѳ����c*�sɈ��D�+�r���Fq���WS���aU�M#�U6ߴj[��M�R�6����+*��nb�4;S�p 7%3�\�u:��sN�2�����Z�[w��e��g�ݜ��'�� ���[���o�u����ʸ���}����h��޷�Ȟ[Z^�^6|�&a�j���<|��h��f�"��x<8�2A�XSpq�D���oK�����8�SU�,�,���G��+!��x �m�/�;�@Bt��%�Q]t�&�n�Ť��������f�0���
wh��+�<W)g�v*��Ae�Ln򩆧h�~Kg͟��F[������ƨ�������h�_������lJ��MT:�V ���BD��E9�U%!��Z�|�N�9�#5���rFN���s�h⾴�J�dv����|�E�VT�
���"MQb������Z�L��Mԅld��*�͘x� �>,�|�*�̚ͅ�8��q�'or	o`]���N4s\���3��l
��/�y�a�C�D����y,���R�Pq�&MO1'�n���>���!r��`Jr�Rևt<b�V<f52�k1�S Y���<ָ���x���W0���1@��������6��l��e��BU=�t c@�r�����Y�)����Vrh�U��s�����+�ӃΓt����V�8������*����NE���YzbqFH�]�'f����&v> Ώ��i#�=��%�7��K����B=0���R���v#m�'����2��hQ>n 88$�g ������>+�N̬dD(��X��\���m�_�,ɪe�6fm�3��Y��Y�e��O$����O�M[ST�6���gb��֍��L$#J6cf�T�e+�B�#����?},1�{�'�02�lQ&��\�Ĵ��/A�(|C�<�O�T��U�i�8�� ��x�?Pb�$;�1?��C��A�B�K�J���K�?͍����y`�O��3g��e/!	���*��mXxo�汤���g�%2���� ����?48��!���hx�esH�jB(��{��#f���SY��,[,̉ZC�Dm�:�j�����3�,����X���JE2M�Z�=�2hc�3S��1_	��@����2�Ȉ���qԦ���?$P�����p⛉<1����Ihz�3��vs1+����������M mK�V�/K{	����\9p��ܺ~p%�I���^I���e7o7����X��5s�+&�UB4�������>�ȕ�j��?�u<)��?�3�6҇Є=��~��Y�Z�n�����ܙf�q�!Q���+�q���2}sĤ�s-��AyQ3��j~���wWE��%�[B��j��|���p$��q�P��
i�<�jUId�YZ�^��+��߶c��,�<X�\���L����v�w
�'~����H��*	?��W������%[��Һu�Z�H����/J.�K�cP��v�'�U��U�\zՕ1~�5R��qM���"(JAI:89��_Shv�kE��ئ�2(�I�CJ�lU�ՙ	�zM��yp�s�	����y��~�d7��,�S>�3�ݱN�7�~�,�S3Ҋ�	�
��Wy�'ǆG	g9L�FTiҍ��icmԭh�ϴ�8�/�r��-)�����T�(xe9^�\�uG�PYK,Sى܍�����%id���'SΥ�ﶞx���N=}�.<���$Ǟp��eAD�S W(?��]���$��ŀ���j(&LG2���"�F��ᒳ�Ե���+3�N��B�?����(dr^B�4�H�@oF�-!��#��$��XE������Z$8�e�T{��O��L���n��.��O�<7�މA/z��7Ni�aU�^���l�o�⎰a0�D@w��1����4������:�e:�vń%#�5w���pv��Y3O�d�M�;ęI����p_����.�Қ���i�N�RPf�%L���z�z|I��oŲ����0��ax���x�U�.��N���8`�= US__UM/�rW��t:�E�0�w_7�u���0K��N�A�Th'x�Lך��Q���n;���=�e0�=J{�"�H{��]=虡����8�kp~��oط��-��^����NU�S��̏ ���
���ς�t}H��ф��I�Y�������������8��^�����#QH��b#�����������gnc���&e�ڲG����]￴��M����Y�?���V�+��2�h��� 2\0��8-j��$R:����@=Z��g�7ǽ����OR˱�؟}�ﭑ݌�Vi�Y|,<S�����Oj`�W����a!B�?$��c\�GϨ~��d�V�I��0H.�wSfR�pW��^�Ve+�b4|��]<]P���P?�r8;ǝR��'춅�dM������>ĥ�u��	��	�$��~ꈏ$�XN?�]�I8����l��&L��m�e�#�g=o�����<�n|�=.G^c{�����8Qᐡg����:c$�e_ݡ��4eH!2K��1s}�qi�D��$ݲ��,ش	b_f�)L��3��Ւ� 3ؕ�ZE4�j����%0�\�(3FW��^�81��25kc^����+*LA%�l��I9иMջݕ���J���s{�GNbd��'-��Q_��5Ub��&E��w$'{I�\F<}�{�Q3w܍g:��e{k�V�dA(� ����T)��D0���ө�~��U��L�#Fp������9R�T�j�0������0���˥�����{j.Xos��jG�Y�k��1B2����O�*˲�h������� �lՎ��+C�ۉf�@���2R?�4>h��AE��`�Z�b���6Yۧ33`�K��}�&�N�jB�
<���@6vsk5��%���R�ң����n���-꣝�si��穳C*�َ��"����.���4y6���m0��gM�0)[�W1��hF���C����5-ƝV4�Nn,�0�W�gٲ('é��G�R�*���uI.'������*;�y~'7��N�4�Ns���qMw����3�!Ӷy�)�崶
�N��eo�m�7�m��}��D�������o��O�N!4�aqu�Xu�bw���&���'\��6�ZJ�ִ_�m%x/W�T�J4�[���ӣ9�[�c~ê���GHv��~�)�x�&�|��
Q��
91=����z��~h4K�]�r�S�5�j&���h��+�%㞣��bX�����==?@���T�#�\�Ix7��������y8����9B{btHP�2����g�j麼�^S��&�ߢ�=�����N�1'C���"�j�H�)~u-�{�(-{��Z9��2Qf���ӽ��.���°��<Iq:a	������]�ϧc�"$��
�V�t����ļMMG�!�x<*�
���샛���X�#j���'Y��g���@]���X��*g�ʴM��ۑRrӎ�~s���j�ra��k\17>3Ԣ�rj�C��&X��'��_78t����*�:��$ǶO[~6��2X���0p�~?��y���)�1��TR�+��v)? 	h�ʫ'%j�7�.^��G<4s���=��[�C��Í�hR^�"�=0y��e����HE6�C���-@ϲ�`��!7��:�jT���N�b�㭵���Eg�\v���K�Xxwr��X\QS��w��0G.Y�{%@��|�w?�w�Q��.<^p��l���"i�4�ZvH���Aǭ�T�Լ�2������ߦpx�;���!#,����BV�n6"x���^=���֤����0�tY���X�[A��M[��v{;}7��[��M�n� l2g����ŔA<�V�����JY�*���+6S�J��dd�h�/l�]an�˰¿�Sø���R㼺Ϋ�tɲ��s UN�nT�6���X�9}[n�ul�2�V^��8���D�x��v`Η�ҹ����a���T�LMW<�yT���'&�A�Ң,������Ő����<Q���Y�w�7Y�s}�o+� ��OIO�K�Q�RF�7F�`� k�|e0>��v��Ӧ���N�EH�J��-Z�fa@X��B��W�t烹(�V��,W�V�/m����#�𥃢�X��Q�=7�k{0�7ދ��3���/��]�﫶z *ܫ��t�t������_iۤw�V*"��x�vb5��mL�Ya�i�8H�1$���ݹ��K��w�StCڦ�VZ�y)��j�'���B�r�w')ME|@ 3N �{e����o������i�nK葨���:uE3����41c�jP�|��~� E���2w�h�M���C�T��I:�5��Ƭ��k����o�O9�Z����J�	ҰQ��[�\ ��DBy���h��OY/W��kg��1�Ā2g�����[��q��t�����4��u��,�b�uznFS��Ĺ	����?Y��?���A4��s�Bq�~7+F�f��_�VE॔j��?g��C�R�?��\YްP��U�*����h_��\j�^;!�����!M}H����y4�\��[�A;-�����nBEY���kfG�6�������r�N3���s|5ݝ�cn����Nw)ߊ��ms��ЙEv��GN==I5��b��۟ʰ��&�
	��o�怬 钃CSr��iU���_�v��>�a\�[8������㶷�Z!L�.��5r٪��8W����������*n(���)\����������u��k�yn����k�9��х�pf�YkXr�*z.��t`�]jKh��a32Rqe�*d 3����?����0Y�����odT�MU7p�Hݦ�s��
;�9�u�������Imϩ[ͬ��"�9Y�Cm�t�`�KT�1)L2�f�)�훝ԫ06�X����`Cp�F�SM�Yc\ڽ�4�+UWV� zi�.uh����66�cU���Q���N,�x�����u嶂�T�o��j
H�VA����=��e��33��g�S�C�b�P���A�QU%^)������r!>E�������ޝ@9c�iT��1|�*{�!?j����}Ν��GӢ� Cî� ��ͦ�E&s��_T��nJ� ٫����S7��fRR�����ݳ�_��I��K�@������{�_�޳!�B«��ƧGA���Cȿ�3��e

	����r`BA���uߎ#��S�| f�jg�jjf�f�g�>�����o,�������g��)S>S9S��pu:��S��i#ȭo��f��hDu��C5����Ro�����w��r6�S�}2���}�c���e�:O���Ĵ�t~�9�`�r�v+�f���x�J� d3o��co�=��<J呥�_UKSE��O���V)��Z�B�#_���;B��`�k0�g��@"�Řg7a¡����D{�Δ�������x�醪X��f8[��AᎥ�����R��\�A� o���6E�}:�J_��!߰.D��.��'A������TQӗS@M���l�_��;u�.��Jm#�����g*�'�F��5j��i����ȷ,.���ǋ\A�`3���n"�����^�`4ذ�%e ��9��q�x=�����5��DšÞ�L�3fC���h�λT%Öj�=a�IT��rL�S��J��kˈ`�m6:�c���!I9�s6:F"�V�%�~�)h�ud<.	g��5B��a檥W>&hx��VU���w�C/+���H�r-)�j��=5�/���]]���a��=��ef(��ߑ���E��5����z���ܢ�QPα+��Y�.���$,E��@;���L!�o�[�|}�U;��D,�w3.9�tSF27d.�f�#5,���<�޸�W�f�EdD��^᠃�Խi�v�f����fX������(HV�Gw`�]t�����$\���"ҕM>O���{Y��kv�s)�Yzv�.���V��͂/�����y�S#���0� *i`J�`? �|���L�O�c_����q�@���^ K�i,��S�P:��CCw\��)F!P6���qwzd6ɨs��_wg��#��֋J�<�:�.H�+�d�^J�l�E0��/�T;�i2`'�턬�\��ts������\�m��8p��J��	g���}F,,�	JC�Kd��-�)�8w�w��>DW��!M�p��F �~|Y�a�+��	?�j)�U�GL�{�<@9����sfDJ�j���C!D��6jT�pw��\��u��2ǟ�q*w�b��0��9Xnr�'��TV�i��ۺ�$�#!̙���tc�d?�%a]>:�sÂ�ۇ�����2@��.v�1�JM���H����W����r�l0���<�+v�!#2"��Z����{��[e\�%���%#�!Oc�(A-3`��\+��6=���XsM���&�%$*�.�
�W�}�ۊ����D���jt�0M�7��S���eL��]\�*���A10ve��'��j+��L�,�s�LwH��9_$��5��G�XH�j]5&�p |I�`4����b�t�Y�_J��}73�o���L�&M������#�|�$�"�i��KV���cdb��oBl�L+=�K��y�aN�O��dCu����t�t�@�j��N�v����M�A�f�����;�|�E9�TBHi�VS�m�܌D�Q�(�zr@;'�*bĈ���D� 7���B�)\�B�R�O"<jC.a�kJ/P~�|�Lg��83f3V������z�v�U�y�H�Ko�a��\�ǏcoY<�e=�����G�C��u�z�=�o��p�zUhB{ ��\�W�Vb<�匙&!��Y"݁o+��յԧt�桳���f:����PT����AY�
�mI�5�V�qB��G+
A> ��6�b���Ҟ���j�_9~J72�E6<x�]omo�$��������bb�jQ&��7:3kNC C��c��'�^$�0�'L����4�R��[�B_A&�0���6Ay�Q�m���8�.�4�z��:�iJk�A-��5�o�}��W ��W��k��#����:.�G7��SXο���E��I	L�`�m�����Q���Bnm�wT��?gx-V�
�r{$��m�ٜ�B�c�63P6���z4�V�ɶ ��ӭ�Lh̰��e�H0�M�e�}��Y�4�[�)��HU[3i�$6�*��C�@H7���]qѻ^q�f��n(1����t�
�և)��Ix�3G��#���7���(��N\%���&�|�٠� ��UjJ%E�kC�8z��QY���o�%��wkTQ �03�A�l֋�G���v�\��M�1����P0s{��g��C�������d�6�x����h�m��@LR���>]Ë�!�/��6�_+��?hBTLle�k�y�Ҵ��|W�@�=�*��N6Vu(�ڀ�gZY����(�R�%3U�:���G�0z%7L��ledv��=���J��!(����B��_㖋�'	�bA�#�/!}����4�25]"��p��KZq�G o��� �p������
隌v�]�5�4؉�ߧ�l�%l-W�eU��@VT��'�ph1&�A�atO�:��ĺ�xWT<.J\&-��������2r�hr�J��<����N�8�!�'���R�*gּ����\MU���i�N^��e�FHAjJC7������[֐���,�7-�l�j7�ԏ�E�����mTzL{r�K�>�:�����ݛo�aB�:��ٍ� S0);y�d�u�!��+��wU�Tk[���m��a����b
�V�ҭw�������29w�6x�"a?���o>�u ��j�4��0�_�n]c���O�&m��3�\�#5��a�7�a)Kh�+��=�i��চ!���Er&K��VA�
H�"V�өP��b�=�9��h�l(��K�D�3W���+NV0Kl����9��\��`	�m4���Y6��N�SnDa�"�t���C`L5����@�3��T�0Y#���^��e�P[�<�krP����� �1�pj�>�1c��o֓�3��&�&��O �s����X|�[�/�"�5�H�5~�kg`�=�� �<�E���`;�T1�{yP�o3��u_��g�<Z3�]S'��{�d1�M�Vk��z�]�%�È���ĥ��� Ec�s=��P�;c6y�]�e�MGi���4�� ��ڧJ:�N�*��|�Q���ŦA7��J�@�7������8�����?�?��c]�p��<浿)l�]�=�-����U���/�����S���%��j��;g?�/��R�|i{�������?��:|� ���!v�_+��?ݞ�(�Ӵᖫ��Ϣ��@/�E��K�O��P�[���"t��j����`��g��U�\�m��ϢU�녑�dh�П�T�cSA�T�'!x-�S��Q=���#ǵ�JU�;�g����N��џ!���9�S��3���O	��-��vH}��w�|Vr�m���}LOO��R!���ijL>m4���������~�
�5 �WF�T��~�Lƿ}\=u�;Hi`�����aD9�F9��>e���������[qla.G��믦b8��#8J��c����Ź�g�^����[@�멢|N0п�������j����X�G�Xp=�s����~���(�_Gp�c?.�)�y�B6]�����(��(Y�y��Ƹ��������Ȧ��t♆��qũ�>���;����<T�y1�"���@�R�b]�#O5��K��p�~^B���xy]Xޣ��=�.���%��;6)Є� #3����o�4g��I��-�m�i�%H㖶�n�b\hE߅E���l�@@��Y�+�����5,�R�  ��((���)�OO��&��B�Cl~׌(oO$�g�D����C�����fj��y|�������,9mT1�$8A+6��q��(�s\/ߦ��ckmH����W��Mׯ)C�L�T�����z�E9q�
��ە�������2hcړJ6���OKn�P��E�wh���E��Y�ʿ���T� �~,S�B�b�%��Jֺ���`ގ/����i6��_�Ti@
x�ۊ�`L�����f!A�@Z�7e���<x~��Yc��p����ު���%�g��)��P#�sS�%!��WI	��}�O:ňU�j��}.��1�]7ͻS����fo�<J�-oD�0bP���&��b6�������"?3�D ��x���d�p�D��%��Q��Q[�d�*����"J�$yk�&
�*棽� �l��u�m��]X�fy�/O@i��!y���,�b��{
�I��@n �%o���k�K��"�/Dl�Yb]៣��� X*��e!pX�f,�Q{}�I#�9.MY �)1�4X��$�R"�wB��\b���K�:�>�b�-ºt9�s|v:3�&��oV�.
yV?�aU���|���;u�{c���x�����Ej.��� �$��AWS�����Fs�XX(BW=,�ݟoC�w�l�'�C�/h|d��|��L-+c��/?�DXu�'�� �FMҾml!ïw�`l{#��R�l�j̬��YL����Q[�W��9!�5	4���szO<k��9�X��ql�=AC�S��B�y��-�����;��/;����k��{��}ު@�ק��|o�<o�!i{r�
������7��P�_����l'�|�c^��	�dʔ�G_�f]&F�u3"+���-�i4�k�:�Io�����z�n�C�Al!ͷp��B*2*�����]S Q:��������kK�g^j�q�)�a"r���vԻ��U $�h���൜�F`��� �����
ٵy>�=Ȭ6�t�.3�� Y��[`�s���->�>y�Y�s� #����Kʅ뫨����$�x��ËA��0�	G@DPPv�zQ��r�W�$��:��ທT"���� ��P38�D�`E����� h�8��v���Yܭ����6�ѡ�[�����u_d\��yO��Ւ�~Ѕ�\_����x��C���P�L�����)���	���x��:;X�]8W���OSߙ��� �I1S�62{]�~�a:���6��T(���2�&�I���F"�X�m�㾵�rcn��/ ��#"��,��^��R��	|�������!7�E��+�&�X]����k�$�Hݡ��|��Pj�T�
�H�EXJd%�����Wi=R23���h#M�f�g]x��7cݶ�L�A�U�҂#Z�s�2�	2���L@���S0�*���n�d����kk;��4��c�T1��B����I:M�y�M�ҥeІ��rrv麝�s-Ev#̿h�ٜ����_��6q�Z����k׍�A�נ�݆�¤�:�d02���B��Q�A0�����vY��s��?Y��RB%֐/�40����\{�|�`iH��]��ȯ;�8QE0y��\���v-q.��׳��s#�hU��h��&b^�(�׳�޺9�;�B ������=��g/�\@�B��9�P��7YNx[v���^�;ZA-2�����ږR8z�~Ä�Mq�vk�X��y�,��I+�MO}��o��J0�u�B��ڭ1y.�Z�L�J3^7��Z�$��҉�p�RUϕ1z./a����Lʝ��i�=�@�Q�a	�|z�,{L��>���� �������3od#ƿ��5�NB�͜�4~Z��lɇe����\ɇ*�f��c�ZT�e���.��L�_��_yj�0A,��!�V&W���u!���(��͢.��,���Ob)oxgJ�F=D��}=�H�Y�f98��Ż��@t������N�n	~�V~|��/Y��; ;�x,�ߓ:��8�|�����~�����-��V�'����fYz��sH$�KktO-�v�Kh��y�
R,hZ��r��
F�P�
��MAm���d����چu�%�6��b�u�C&�cs�-������G�m�-!��嗿�#L��t3I�jM.s��[���a.&�-�wr��5x�0�~{���e>P�b�d��(<��5!{�-=�`�
��*��,=30�Cڌ8��A��J#n�"����8`�{�NU?�Pt���>*6��W4a�p�����k��(��GVr���S^r0���3$OVyMj*i��wȑ�h�82d\�*yvm�w����	��������5���;Q��*k���U/B�t|��X�dewm� !]`�m��H2����b�{�"
**�~$kxUc�HGʭ:5���X���9<-�&�G��yb�*��X~,m>qTcA��G! 4�l�j�L1�&���*ۋ��Pj��94M���6���ci�X2�ER�[5��n`�Q,nY��iAj��_��w���YA=P�&
�HH,<L��Xf��bw���M �01(�)!c�L[����&\�����8�4�
��_[ۍ���i��^&C��	��
s(�����1�Xݮ4h�ql,�
��)CA��\�"��-ix*�8�*1k ���P�	V�\M0�����L���5b��n����[?�
Ї�������ߦn�K����E���K�FUC�"2�c�B숩�P���4�
��zQt�!z�������\�Y��=#lvAk �`�JCH�m�jz��N��P"�)f�`1�ݱ� �c*?q�%��@��G#���r�v��s� ���!㚃�xhB2Y��U�T��f��WR�Ii�SԨPN]�T�W�nM&Vy=�-d5�(����J�l�Ƨ1{W�K��
��=�-�Z��5�K�@k�H&b(�,�%�Ʈ�� ����a���TƘ���l6��|DV�b�#|�\s�߼#�H.�v��:��x�2�Z7���Q����/�2����3��#����觮�����)�g.k���Q��s5�*�p���t� ?�2�����1=��y�����o2.X�ߴh����j�(ea�5b�/�Mn����k�(ܽ$I�	C=�>\{�v�}���1+\ �U�d����K��pv��B����o�̐�C1K�"�q�NZ�KH����^�#��DD���Ƚ� �*%�# ��D%==s�[B-�f�F����ƞ� ��^<�fV�j��A����h�ץ@׼sV�/�Cv�W�8!V=%��*�K�kn2��"�/�b���aG)d�d��3��Q����gY��1J���}&M(�N�A��{�h3-�Y|��R���V�z�|�r?�&�Ľ61� �C�i��9;b1���	W�4��~�=� �_�A��n^�A��H��U��M���D��Z���`aUx�����x�BTo̪�R�f�=�"��Q� ����Գd�E�+��4S]�gҥ"�H�V+j�� �R���~����)�?r���)�?r���	_��� ��� (      !1AQaq����0�����p��  ?� � ȝ�1G��������?��S���?��{����/y������ �O��������� �?��?r� s���?T� r<���Z��N?k�~�������=���C������/��!��{�޿���f%]7;1ߗr@��6	�n�b�B&6��XC.�;���z9�9^�ӓ�X� S7��� �nY�x��N�P��ĕ�Z(|f������W�d]k��Ez��}L�����4M7'��::<�8P�i8 ���[��m��_:�sf9)$� � �M�̫�|�)�kWA�Iyp�&���l�E|�ph:S�<ⷤI���$��Ke.#���J�!�aq@S�`.+�׈�gxjKp�y嗬�W��=q�Z�O��8C�5��gy��}qi{���Nqr�����]�黟6I9S��e����]����W.E�E�¥��v�S�:n*E�:�LT"D���	���������띊�F�Y v��S�p|c�0�'�A����=�����C�@
6��0�����PFn���g4���(pf��������g��!+�"]��&��=vg�L0 W.y.�c xk�W�ޭ�(ky\ �YT3��{�K�k��}x��Q�?�?C��T<b���7�c�d��!��MI��`n�XG~����c�x܄m�S���6��Ć�,y��^n����]AZo�Dުe���'�}��/Y���ԲDK�xwp��8V���H�[�*��8��5�����@,�������O�6:��D|��0#��� XI����t��!�S��$� }n]��E~"1�(� ]�Ď��b�B��-�`5�U��r�3˃W ReL7Sض���$���<��\
�����:�9� �
ɰ�!:�+��E{�aV������p9Էo����#����]#�f[�H�:]99/8�_xd����� �?Tb
o��w��� Kш�+}h��:�d6�-�Ʊ�X���i5180&��k� ��"Q��?�~�`�?\� � L�`����c���j�H����G�i� X�s9����=�q�.��KxY|"c@oXG�n������F��a}�3�o���� �'�~/�?�ڡ�N�
5%}��@��G����6�Z���#�Co���`$��\To9|騬!ϴ���c�/8  �%cӓL�p	_Z��_&��Ɛ�\c:Z�I�8�8�.T��y��� �90T��TP)>Y�x;��
��G��c�ʻ��s��tX� ��4C�9Ɇ�[?��,[c������H��]`�H�F�� s-X�c�Zv����S��w5��x䅇.�4�����5������u�r&�#�n�=��
#�f��TGk�),-�L����:����dw��y��m�bR0�&�N[�in�)a�2�D�1�� yX��L��3@�I �x\���?���_����yʃgX��@��(���@#mʗ쁍m���7N���O�����w5�;��� 2�������^��+���9�`Z�VbR���y�	�?��Yy��o���<ܦ�\32`��|�<D���~�~���J�`��e�Ŝ���� y� >��t}�U{^� ����z�'��X�s�9yV�G�� �Y�G�����%�#l�h^�� �/=��f�,5�_���+�n 5��9�|ʋ�m�?]�Z(%d�]}��U�}�"�P�)�~1�����h�!��\�a,G����+:�Nkxu������%+�N��j)�i�1���h���Zw�r�� ��=f�uHGbr�h�n(�C�&��� *��"� X�a{8p@�  mۚ��g���5��[4]}p��M�}� z���4�Z�nC��Y0h� �G\ky����J�p�I�(J��M_1+�
�a��U�W�����6�#c@`�Aϒ~&)���9K�U�AZ:�7i=M��=cW. ��7���\���^�q��u���R�$^�"��;Zx�#2�X�_�[K���G�7�lJ��@�Ӄ��n����B����}p�R_ z|�.��P���ƨ?�b+xT�I�L���n�c�E�FP+�B9ް��d� ���@b-�ޠ�����œ���`p�A�Iȁ��:�vN�i�p�cwI���	��(�s�`��7��O��a5.�O��8=�l�Ŷz���7�{�.HO� pBO/��%J���}0��T�cF�n������y����8)g�)@�P)8\m��ʍO�˚��0��ȀX�o&^qQ]�&� ��z��԰oj�׬��Y�C�dd�`vT� ���sD�o�*��{spV�(��p����z��s�Z$o�Q�J���d�u�h���/-8��"���|џ�=`>��I@��0�U���rOd�/��Q��+az�t�kX&tM���)�F������O�D�j84�t�X����]&���{� |d��L��%�z�50�7�e~����۞�~���t��x���j��,>�L�爏���W� H� X4i�I�{a�R��#�������3I��G���xx���M~� �(��M����Į��+\�@Ȼ��>���	t/�܂C@���p7@I�������������a��-~ޱ��7���ë1O@�i\@�+���`V��vb�܄�O��1�	d�vS�XtQ7H	�ޥ�ID�ԓ��Gx:l����D��W�I��#��x�H�<38�<F��!�|�Z�p�ѝLjO�_���&��	��Y{�6��:��Ϝ��Z����Ji�H��{�I���lW'��� ��2�{�_���E�"��0��μ�*wv]۳��%� 8U�w��OT�\�K^Y>�42X)	�Q�hrC�bo����f)��豱�	�7�W V0��>����*��n�'44e���'�����:�:N���=� �F/R��K��� �!���:{�4!�@?Ɇ�q�#x�>�Y ��^�ظ�F`Q�وĂa k~\D�$�}�<"d�����㞱�r��^�pY�S�w�~�F
��>�`��(M�q;Đ ��=a���RJs&j0Yp��7�>F2��7 (�]":��  P���־��k���4��W#0D��]��x -x	��� �\�� ����N�����8�Q�Z>�`�",O�-8���[�l�d�Q�������Jf�bw�Y�j.Ny�N��>���3�9+�Ǖu�j�i�x�D碎�.Vrȉ}�4v��+�|vb�8\W���gV�Ԥ�4ݤM�G�)�T�]�eO�)��6���k+�˲�� '�j��"#��OX����%h�ϦJ@Z����$��	'8y}�l�M�A�J���-��I)�}L�c��U{�^�y�Ӻ\��(@E��|L������29�������vx�"Ճ�p{qǇ[@��p���Uܡ�ql���	ъ��P�4�ͭ��O2m>LMq��6��ȼ2@*�?8�9���*��!�7L Oo9��)Xh�a=ʝD N� #уFkK��
D��h
��D%�W������z�zǢ�0�]�(��'���Z ��o|�u��$t��~�.L?��?���C��؊#D�ĚP8K���H� <����G$SM M'fm��y'bk&C*�[���lDy8;r�����I��!�$�y�0іb畐"1_I��
�>7�A����w���-�m�Z=� x����4��/o�9���H�2	�8�����u��Wx,�U	����?�Ï����8*R_Vď-3!d��4n9P�*���RQ����9|],����'�p=C}�O�&q��>���� �X��7j��ϖ��0��½�����چJb�·�4�h(4na5P6r}z� ���`\�	��d��M�^q�mh�x�dTbة�&�l�$�lm�4.a>�̊j�ҥS��	�CX����EK�*�Obq$��XD�����\hO9CD �\�]��wǬ���E���4�����yy�H�G��v�#Q����&ŭ�C��I\D$:S�9p6�Dy5������D�{77$	D:���M(���f�dr����o��Ȓ���G�F��G��56�6��|9ʨ֝���v��/���:�O�bvf�CkED�Bf���lr�e�(i�E�k�a��_��|���п�1��LHH����a&���H7`LT^8)����r���4BaUX5ǚ{�E�C���N�PG#����,I
�]F<R�����0@��7�׼"�Ǥق.��8�Km�W%]�ߌes�A���$�QLO���h�g�ƕ��(�瑅���a{&���(5NGF���
CH��Kܓ�7�L_�B����o�p����u��Z�|x�0a�h��yņ�ꢅ���/�S�깈�������A�B���j��[��x(Cs�_L11Z%EO��ZA�@�.Q7�S?��=�!3j��t��w�z@��Y�8
�q��p�T�5	��$}bA��
�:o�oo2@ó��@�� tF�:�-A�T�^M{��R0Z��o%=���tw�9�t(��zñD�.��5:.*r=�gN̰^�S�`.��m�A�펪m��?�����n�U����Rf jqw�-��y��Nw��M�~P%T|����K�� !�� �5��~�����?��~׼�+��O������?�y���y��>�������bҟ#��{��`_e�/��m��=�Ӂ���q�� �_��PK   c��TXK8�  �     jsons/user_defined.json��Ao� ��J��F��6�M˥�MS���hr0���nE��{N��mZשw����xz�v��6�Q��U��X]�=h�� �`
;�[�G��ܝ_��!����dZ�4��֮u~Vz�pX�]���V�;� ����n[FȔ�QBU�2De1�i�9Kc.� Rh��8}���y�;�X�B�M�?��ͨ�x��{�k����C���zaBS�Ϯ��#ʱ�,'p��u�1@[�Y��My�z|�i��W��԰�p�%%�D�8��n�'�~;駷��J�h��Cp��*�0���r*<��S������>�.�蓻��'7&�gS�� |��8��DL��˿T|��<���Ѳ��Z{��Lٚ�O{*g��T_�s7nZ]�Kw�q�ˌ���d�ƼȊ8_�p+g��sJ����1��"#\�j�s�J�r�q��,�X"0���(�3�����o���T��p��>�~팏��r�PK
   c��T�t��`  �                  cirkitFile.jsonPK
   ���T7�I� �" /             �`  images/39ed726b-0701-4a7a-8bd7-442054548109.pngPK
   &��T��beY  �[  /             n images/c5cf112c-a0c7-416d-8826-4525095e4ef3.pngPK
   c��TXK8�  �               �� jsons/user_defined.jsonPK      <  ��   